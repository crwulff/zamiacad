library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_misc.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;

-- This is a small hardware configuration circuit which also contains
-- other misc stuff that is not worth to build a own core.

-- It allows to set or clear a signal to configure the Hardware, e.g.
-- debug_mode of the switch or to set and clear leds.

-- Also interrupts will be controlled by this component.
-- A simple timer is also available.

entity hw_ctrl is
  port(
    --generic
    clk : in std_logic;
    res : in std_logic;

    --io_ports
    hw_ctrl_enable : in  std_logic;
    hw_ctrl_dir    : in  std_logic;
    hw_ctrl_adr    : in  std_logic_vector (13 downto 0);
    hw_ctrl_write  : in  std_logic_vector (31 downto 0);
    hw_ctrl_read   : out std_logic_vector (31 downto 0);
    hw_ctrl_ready  : out std_logic;

    --leds and other misc signals
    hw_ctrl_leds        : out std_logic_vector (30 downto 0);
    hw_ctrl_ledl_enable : out std_logic;
    hw_ctrl_ledr_enable : out std_logic;
    hw_ctrl_ledb_enable : out std_logic;
    debug_mode          : out std_logic;
    
    --outgoing irq_signals (to cpu)
    irq_adr : out std_logic_vector (31 downto 0);
    irq     : out std_logic;

    -- input for interrupts possibly generated by HASE
    irq_input_softirqs_com     : in std_logic_vector (30 downto 27);
    irq_input_softirqs_pcdebug : in std_logic_vector (30 downto 27);
    --incoming irq lines
    vga_vblank_irq             : in std_logic;

    --buttons
    BOARD_BUTTON : in std_logic_vector (2 downto 0)
    );
end;

architecture behavioral of hw_ctrl is
  type states is ( idle, reading, writing);
  signal state : states;

  subtype mask_type is std_logic_vector(30 downto 0);

  signal leds      : mask_type;
  signal ctrl0     : mask_type;
  signal mask      : mask_type;
  signal read_data : std_logic_vector (31 downto 0);

  signal button_old    : std_logic_vector(2 downto 0);
  signal button_change : std_logic_vector (2 downto 0);

  signal irq_en       : mask_type;
  signal irq_ctrl     : mask_type;
  signal irq_hdl_adr  : std_logic_vector(31 downto 0);
  signal irq_activate : mask_type;

  signal   TIMER            : std_logic_vector(31 downto 0);
  signal   TIMER_RELOAD     : std_logic_vector(31 downto 0);
  signal   TIMER_DIV        : std_logic_vector(4 downto 0);
  constant TIMER_DIV_RELOAD : std_logic_vector(4 downto 0) := "11000";  -- 24
  signal   TIMER_IRQ        : std_logic;

  subtype io_adr_type is std_logic_vector(3 downto 0);

  --mask adrs
  constant adr_hw_ctrl_leds  : io_adr_type := "0000";
  constant adr_hw_ctrl_ctrl0 : io_adr_type := "0001";
  constant adr_irq_en        : io_adr_type := "0010";
  constant adr_irq_ctrl      : io_adr_type := "0011";
  --other adrs
  constant adr_irq_adr       : io_adr_type := "1111";
  constant adr_timer         : io_adr_type := "1110";
  constant adr_timer_reload  : io_adr_type := "1101";

  --bit to select pcdebug or com mode    - in ctrl0
  constant pcdebug_com_select_bit : integer := 0;

begin

  --mapping of irq activating signals
  irq_activate(0)             <= TIMER_IRQ;
  irq_activate(1)             <= vga_vblank_irq;
  irq_activate(4 downto 2)    <= button_change;
  irq_activate (30 downto 27) <= irq_input_softirqs_pcdebug when (ctrl0(pcdebug_com_select_bit) = '1') else irq_input_softirqs_com;

  process(clk)
  begin
    if clk'event and clk = '1' then

      if res = '1' then
        state        <= idle;
        leds         <= (others => '0');
        ctrl0        <= (others => '0');
        irq_en       <= (others => '0');
        irq_ctrl     <= (others => '0');
        irq_hdl_adr  <= (others => '0');
        TIMER        <= (others => '0');
        TIMER_RELOAD <= (others => '0');
        TIMER_DIV    <= TIMER_DIV_RELOAD;

      else
        --timer
        TIMER_DIV   <= TIMER_DIV - 1;
        if TIMER_DIV = 0 then
          TIMER_DIV <= TIMER_DIV_RELOAD;
          TIMER     <= TIMER - 1;
          if TIMER = 0 then
            TIMER   <= TIMER_RELOAD;
          end if;
        end if;
        
        --compute state
        case state is
          when idle =>
            if hw_ctrl_enable = '1' then
              if hw_ctrl_dir = '1' then
                state <= writing;

                case hw_ctrl_adr(3 downto 0) is
                  when adr_hw_ctrl_leds  => leds         <= mask;
                  when adr_hw_ctrl_ctrl0 => ctrl0        <= mask;
                  when adr_irq_en        => irq_en       <= mask;
                  when adr_irq_ctrl      => irq_ctrl     <= mask;
                  when adr_irq_adr       => irq_hdl_adr  <= hw_ctrl_write;
                  when adr_timer         => TIMER        <= hw_ctrl_write;
                  when adr_timer_reload  => TIMER_RELOAD <= hw_ctrl_write;
                  when others            => null;
                end case;

              else
                state <= reading;
              end if;
            end if;

          when writing =>
            if hw_ctrl_enable = '0' then
              state <= idle;
            end if;

          when reading =>
            if hw_ctrl_enable = '0' then
              state <= idle;
            end if;

          when others => null;
        end case;

        --trigger irqs
        for i in 0 to 30 loop
          if irq_activate(i) = '1' and irq_en(i) = '1' then
            irq_ctrl(i) <= '1';
          end if;
        end loop;

        --update button_old
        button_old        <= BOARD_BUTTON;
        ctrl0(6 downto 4) <= BOARD_BUTTON;

        --sync output
        hw_ctrl_read <= read_data;        
      end if;
    end if;
  end process;

  --process for triggering irq
  process(irq_ctrl, irq_en)
  begin
    irq     <= '0';
    for i in 0 to 30 loop
      if irq_ctrl(i) = '1' and irq_en(i) = '1' then
        irq <= '1';
      end if;
    end loop;  -- i
  end process;

  --process for calculating BUTTON changes
  process(button_old, BOARD_BUTTON)
  begin
    for i in 0 to 2 loop
      if button_old ( i ) /= BOARD_BUTTON ( i ) then
        button_change ( i ) <= '1';
      else
        button_change ( i ) <= '0';
      end if;
    end loop;  -- i
  end process;

  --trigger TIMER_IRQ
  process(TIMER)
  begin
    TIMER_IRQ   <= '0';
    if TIMER = 0 then
      TIMER_IRQ <= '1';
    end if;
  end process;

  --process for hw_ctrl_ready
  process(state)
  begin
    hw_ctrl_ready     <= '-';
    case state is
      when idle    =>
        hw_ctrl_ready <= '0';
      when writing =>
        hw_ctrl_ready <= '1';
      when reading =>
        hw_ctrl_ready <= '1';
      when others  => null;
    end case;
  end process;

  --process for reading
  process(clk,
          hw_ctrl_adr(3),
          hw_ctrl_adr(2),
          hw_ctrl_adr(1),
          hw_ctrl_adr(0),
          leds, ctrl0, irq_en, irq_ctrl, irq_hdl_adr, TIMER, TIMER_RELOAD)
  begin
    read_data <= (others => '0');

    case hw_ctrl_adr(3 downto 0) is
      when adr_hw_ctrl_leds  => read_data (30 downto 0) <= leds;
      when adr_hw_ctrl_ctrl0 => read_data (30 downto 0) <= ctrl0;
      when adr_irq_en        => read_data (30 downto 0) <= irq_en;
      when adr_irq_ctrl      => read_data (30 downto 0) <= irq_ctrl;
      when adr_irq_adr       => read_data               <= irq_hdl_adr;
      when adr_timer         => read_data               <= TIMER;
      when adr_timer_reload  => read_data               <= TIMER_RELOAD;
      when others            => null;
    end case;
  end process;

--compute new mask value
  mask <= (read_data (30 downto 0) and (not hw_ctrl_write(30 downto 0)))
          when (hw_ctrl_write(31) = '0') else
          (read_data (30 downto 0) or hw_ctrl_write(30 downto 0));

  hw_ctrl_leds (30 downto 0) <= leds(30 downto 0);
  debug_mode                 <= ctrl0(0);
  hw_ctrl_ledl_enable        <= ctrl0(1);
  hw_ctrl_ledr_enable        <= ctrl0(2);
  hw_ctrl_ledb_enable        <= ctrl0(3);
  irq_adr                    <= irq_hdl_adr;

end behavioral;
configuration CFG_HW_CTRL_BEHAVIORAL of hw_ctrl is
  for BEHAVIORAL
  end for;
end CFG_HW_CTRL_BEHAVIORAL;
