LIBRARY GRLIB;

use GRLIB.DEVICES.ALL;

entity foo is
end;

architecture rtl of FOO is

begin

end;


