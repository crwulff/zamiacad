library ieee;
use ieee.std_logic_1164.all;

entity ccTest is
  port( a, b : IN bit; z : OUT bit);
end entity ccTest;

architecture RTL of ccTest is 

    CONSTANT decode      : STD_ULOGIC_VECTOR := "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111110111111" ;

begin

end architecture RTL;

