module foo ;

/*
 * longer comment with `PREPROCESSOR macro
 */

parameter dw = 42;

endmodule
