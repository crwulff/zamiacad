module lvalue ;

always @(spr_addr)
   a[5:0] = 0;

endmodule
