library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_1164.all;

library std;
use STD.textio.All;
use work.manikconfig.all;
use work.manikpackage.all;

library UNISIM;
use UNISIM.vcomponents.all;

package maniklattice is

    component SP8KA
        generic(REGMODE    : string  := "NOREG";
                GSR        : string  := "DISABLED";
                WRITEMODE  : string  := "NORMAL";
                RESETMODE  : string  := "ASYNC";
                CSDECODE   : string  := "111";
                DATA_WIDTH : integer := 18;
                INITVAL_00 : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_01 : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_02 : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_03 : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_04 : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_05 : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_06 : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_07 : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_08 : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_09 : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_0A : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_0B : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_0C : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_0D : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_0E : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_0F : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_10 : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_11 : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_12 : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_13 : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_14 : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_15 : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_16 : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_17 : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_18 : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_19 : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_1A : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_1B : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_1C : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_1D : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_1E : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_1F : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000"
                );
        port(CE   : in  STD_ULOGIC; CLK  : in  STD_ULOGIC; WE   : in  STD_ULOGIC;
             CS0  : in  STD_ULOGIC; CS1  : in  STD_ULOGIC; CS2  : in  STD_ULOGIC;
             RST  : in  STD_ULOGIC;
             DI0  : in  STD_ULOGIC; DI1  : in  STD_ULOGIC; DI2  : in  STD_ULOGIC; DI3  : in  STD_ULOGIC;
             DI4  : in  STD_ULOGIC; DI5  : in  STD_ULOGIC; DI6  : in  STD_ULOGIC; DI7  : in  STD_ULOGIC;
             DI8  : in  STD_ULOGIC; DI9  : in  STD_ULOGIC; DI10 : in  STD_ULOGIC; DI11 : in  STD_ULOGIC;
             DI12 : in  STD_ULOGIC; DI13 : in  STD_ULOGIC; DI14 : in  STD_ULOGIC; DI15 : in  STD_ULOGIC;
             DI16 : in  STD_ULOGIC; DI17 : in  STD_ULOGIC;
             AD0  : in  STD_ULOGIC; AD1  : in  STD_ULOGIC; AD2  : in  STD_ULOGIC; AD3  : in  STD_ULOGIC;
             AD4  : in  STD_ULOGIC; AD5  : in  STD_ULOGIC; AD6  : in  STD_ULOGIC; AD7  : in  STD_ULOGIC;
             AD8  : in  STD_ULOGIC; AD9  : in  STD_ULOGIC; AD10 : in  STD_ULOGIC; AD11 : in  STD_ULOGIC;
             AD12 : in  STD_ULOGIC;
             DO0  : out STD_ULOGIC; DO1  : out STD_ULOGIC; DO2  : out STD_ULOGIC; DO3  : out STD_ULOGIC;
             DO4  : out STD_ULOGIC; DO5  : out STD_ULOGIC; DO6  : out STD_ULOGIC; DO7  : out STD_ULOGIC;
             DO8  : out STD_ULOGIC; DO9  : out STD_ULOGIC; DO10 : out STD_ULOGIC; DO11 : out STD_ULOGIC;
             DO12 : out STD_ULOGIC; DO13 : out STD_ULOGIC; DO14 : out STD_ULOGIC; DO15 : out STD_ULOGIC;
             DO16 : out STD_ULOGIC; DO17 : out STD_ULOGIC);
    end component;

    component DP8KA
        generic(REGMODE_A    : string  := "NOREG";
                REGMODE_B    : string  := "NOREG";
                GSR          : string  := "DISABLED";
                WRITEMODE_A  : string  := "NORMAL";
                WRITEMODE_B  : string  := "NORMAL";
                RESETMODE    : string  := "ASYNC";
                CSDECODE_A   : string  := "111";
                CSDECODE_B   : string  := "111";
                DATA_WIDTH_A : integer := 18;
                DATA_WIDTH_B : integer := 18;
                INITVAL_00   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_01   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_02   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_03   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_04   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_05   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_06   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_07   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_08   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_09   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_0A   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_0B   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_0C   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_0D   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_0E   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_0F   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_10   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_11   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_12   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_13   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_14   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_15   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_16   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_17   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_18   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_19   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_1A   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_1B   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_1C   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_1D   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_1E   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
                INITVAL_1F   : string  := "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000"
                );
        port(CEA   : in  STD_ULOGIC;
             CLKA  : in  STD_ULOGIC;
             WEA   : in  STD_ULOGIC;
             CSA0  : in  STD_ULOGIC; CSA1  : in  STD_ULOGIC; CSA2  : in  STD_ULOGIC;
             RSTA  : in  STD_ULOGIC;
             CEB   : in  STD_ULOGIC;
             CLKB  : in  STD_ULOGIC;
             WEB   : in  STD_ULOGIC; CSB0  : in  STD_ULOGIC; CSB1  : in  STD_ULOGIC; CSB2  : in  STD_ULOGIC;
             RSTB  : in  STD_ULOGIC;
             DIA0  : in  STD_ULOGIC; DIA1  : in  STD_ULOGIC; DIA2  : in  STD_ULOGIC; DIA3  : in  STD_ULOGIC;
             DIA4  : in  STD_ULOGIC; DIA5  : in  STD_ULOGIC; DIA6  : in  STD_ULOGIC; DIA7  : in  STD_ULOGIC;
             DIA8  : in  STD_ULOGIC; DIA9  : in  STD_ULOGIC; DIA10 : in  STD_ULOGIC; DIA11 : in  STD_ULOGIC;
             DIA12 : in  STD_ULOGIC; DIA13 : in  STD_ULOGIC; DIA14 : in  STD_ULOGIC; DIA15 : in  STD_ULOGIC;
             DIA16 : in  STD_ULOGIC; DIA17 : in  STD_ULOGIC;
             ADA0  : in  STD_ULOGIC; ADA1  : in  STD_ULOGIC; ADA2  : in  STD_ULOGIC; ADA3  : in  STD_ULOGIC;
             ADA4  : in  STD_ULOGIC; ADA5  : in  STD_ULOGIC; ADA6  : in  STD_ULOGIC; ADA7  : in  STD_ULOGIC;
             ADA8  : in  STD_ULOGIC; ADA9  : in  STD_ULOGIC; ADA10 : in  STD_ULOGIC; ADA11 : in  STD_ULOGIC;
             ADA12 : in  STD_ULOGIC;
             DIB0  : in  STD_ULOGIC; DIB1  : in  STD_ULOGIC; DIB2  : in  STD_ULOGIC; DIB3  : in  STD_ULOGIC;
             DIB4  : in  STD_ULOGIC; DIB5  : in  STD_ULOGIC; DIB6  : in  STD_ULOGIC; DIB7  : in  STD_ULOGIC;
             DIB8  : in  STD_ULOGIC; DIB9  : in  STD_ULOGIC; DIB10 : in  STD_ULOGIC; DIB11 : in  STD_ULOGIC;
             DIB12 : in  STD_ULOGIC; DIB13 : in  STD_ULOGIC; DIB14 : in  STD_ULOGIC; DIB15 : in  STD_ULOGIC;
             DIB16 : in  STD_ULOGIC; DIB17 : in  STD_ULOGIC;
             ADB0  : in  STD_ULOGIC; ADB1  : in  STD_ULOGIC; ADB2  : in  STD_ULOGIC; ADB3  : in  STD_ULOGIC;
             ADB4  : in  STD_ULOGIC; ADB5  : in  STD_ULOGIC; ADB6  : in  STD_ULOGIC; ADB7  : in  STD_ULOGIC;
             ADB8  : in  STD_ULOGIC; ADB9  : in  STD_ULOGIC; ADB10 : in  STD_ULOGIC; ADB11 : in  STD_ULOGIC;
             ADB12 : in  STD_ULOGIC;
             DOA0  : out STD_ULOGIC; DOA1  : out STD_ULOGIC; DOA2  : out STD_ULOGIC; DOA3  : out STD_ULOGIC;
             DOA4  : out STD_ULOGIC; DOA5  : out STD_ULOGIC; DOA6  : out STD_ULOGIC; DOA7  : out STD_ULOGIC;
             DOA8  : out STD_ULOGIC; DOA9  : out STD_ULOGIC; DOA10 : out STD_ULOGIC; DOA11 : out STD_ULOGIC;
             DOA12 : out STD_ULOGIC; DOA13 : out STD_ULOGIC; DOA14 : out STD_ULOGIC; DOA15 : out STD_ULOGIC;
             DOA16 : out STD_ULOGIC; DOA17 : out STD_ULOGIC; DOB0  : out STD_ULOGIC; DOB1  : out STD_ULOGIC;
             DOB2  : out STD_ULOGIC; DOB3  : out STD_ULOGIC; DOB4  : out STD_ULOGIC; DOB5  : out STD_ULOGIC;
             DOB6  : out STD_ULOGIC; DOB7  : out STD_ULOGIC; DOB8  : out STD_ULOGIC; DOB9  : out STD_ULOGIC;
             DOB10 : out STD_ULOGIC; DOB11 : out STD_ULOGIC; DOB12 : out STD_ULOGIC; DOB13 : out STD_ULOGIC;
             DOB14 : out STD_ULOGIC; DOB15 : out STD_ULOGIC; DOB16 : out STD_ULOGIC; DOB17 : out STD_ULOGIC);
    end component;

    component latspram_ecp
        generic (MEM_DATA_WIDTH : integer;
                 MEM_ADDR_WIDTH : integer);
        port (clk    : in  std_logic;
              addr   : in  std_logic_vector(MEM_ADDR_WIDTH-1 downto 0);
              data_i : in  std_logic_vector(MEM_DATA_WIDTH-1 downto 0);
              enb    : in  std_logic;
              rst    : in  std_logic;
              we     : in  std_logic;
              data_o : out std_logic_vector(MEM_DATA_WIDTH-1 downto 0));
    end component;
    
    component adsu_ecp
        port (DataA   : in  std_logic_vector(31 downto 0);
              DataB   : in  std_logic_vector(31 downto 0);
              Cin     : in  std_logic;
              Add_Sub : in  std_logic;
              Result  : out std_logic_vector(31 downto 0);
              Cout    : out std_logic);
    end component;

    component ecp_pll
        generic (IN_FREQ_MHZ   : integer;
                 CORE_FREQ_MHZ : integer;
                 CLK_DIVBY     : integer;
                 CLK_MULBY     : integer);
        port (CLK   : in  std_logic;
              RESET : in  std_logic;
              CLKOP : out std_logic;
              LOCK  : out std_logic);
    end component;
    
end maniklattice;
