
entity ccTest is
  port( a, b : IN bit; z : OUT bit);
end entity ccTest;

architecture RTL of ccTest is 

    CONSTANT decode      : bit_vector      := "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111111111111" &
                                              "1111111110111111" ;

begin

end architecture RTL;

