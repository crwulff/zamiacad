library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_textio.all;
use std.textio.all;
use work.mlite_pack.all;

entity mlite2sram is
   port(clk             : in std_logic;
        -- communication pins with mlite cpu
        mem_byte_sel    : in std_logic_vector(3 downto 0);
        mem_write       : in std_logic;
        mem_address     : in std_logic_vector(31 downto 0);
        mem_data_w      : in std_logic_vector(31 downto 0);
        mem_data_r      : out std_logic_vector(31 downto 0);
	mem_pause       : out std_logic;
	-- communication pins with SRAM on xsv300 board
	sram_we_hi      : out std_logic;
	sram_we_lo      : out std_logic;
	sram_ce_hi      : out std_logic;
	sram_ce_lo      : out std_logic;
	sram_oe_hi      : out std_logic;
	sram_oe_lo      : out std_logic;
	sram_address_hi : out std_logic_vector(18 downto 0);
	sram_address_lo : out std_logic_vector(18 downto 0);
	sram_data_hi    : inout std_logic_vector(15 downto 0);
	sram_data_lo    : inout std_logic_vector(15 downto 0));
end; --entity ram

architecture logic of mlite2sram is

   signal data   : std_logic_vector (31 downto 0); -- prefeched data from sram
   signal output : std_logic_vector (31 downto 0); -- data sent to memory bus

   type STATE_TYPE is (
      READ,
      WRITE
   );

   signal state, next_state : STATE_TYPE;

begin

   set_state: process(clk) --, state, next_state)
   begin
      if clk'event and clk = '1' then
         state <= next_state;
      end if;
   end process;

   work: process(state, mem_byte_sel, mem_write, mem_address, mem_data_w,
                 sram_data_lo, sram_data_hi, data)
   begin
      -- set defaults
      sram_address_hi <= mem_address(18 downto 2) & "00"; -- ram is accessed by word only
      sram_address_lo <= mem_address(18 downto 2) & "00"; -- hence 0002 would be illegal
      sram_ce_hi      <= '0'; -- chip enable can be set at all time (ce is active at 0)
      sram_ce_lo      <= '0';
      sram_we_hi      <= '1'; -- don't write
      sram_we_lo      <= '1';
      sram_oe_hi      <= '1'; -- don't read either
      sram_oe_lo      <= '1';
      sram_data_hi    <= "ZZZZZZZZZZZZZZZZ"; -- don't write anything to sram
      sram_data_lo    <= "ZZZZZZZZZZZZZZZZ";
      mem_pause       <= '0'; -- don't pause cpu
      next_state      <= READ;
      output          <= "ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ";

      -- check if this component is supposed to be active
      if mem_address (31 downto 19) = "0000000000000" then

         case state is
            -- always start reading
	    when READ =>
	       -- enable sram output
	       sram_oe_hi <= '0';
	       sram_oe_lo <= '0';
	       
	       -- check if boot memory is read
	       case mem_address(31 downto 2) is
                  -- TIMING TEST - see timing.s
                  --when "000000000000000000000000000000" => output <= "00100100000000100000000000100000";
                  --when "000000000000000000000000000001" => output <= "00111100000000010000000000001000";
                  --when "000000000000000000000000000010" => output <= "00001000000000000000000000000001";
                  --when "000000000000000000000000000011" => output <= "10101100001000100000000000000000";
                  --when "000000000000000000000000000100" => output <= "00000000000000000000000000000000";

                  -- SERIAL WRITE TEST - see output.s
                  --when "000000000000000000000000000000" => output <= "00100100000000100000000000000001";
                  --when "000000000000000000000000000001" => output <= "00111100000000010000000000001000";
                  --when "000000000000000000000000000010" => output <= "10101100001000100000000000000000";
                  --when "000000000000000000000000000011" => output <= "00001000000000000000000000000001";
                  --when "000000000000000000000000000100" => output <= "00100000010000100000000000000001";

                  -- SERIAL READ TEST - see echo.s
                  --when "000000000000000000000000000000" => output <= "00111100000000100000000000001000";
                  --when "000000000000000000000000000001" => output <= "10001100010000100000000000000100";
                  --when "000000000000000000000000000010" => output <= "00111100000000010000000000001000";
                  --when "000000000000000000000000000011" => output <= "00001000000000000000000000000000";
                  --when "000000000000000000000000000100" => output <= "10101100001000100000000000000000";

                  -- MEMORY TEST - see memtest2.s
                  --when "000000000000000000000000000000" => output <= "00100100000000100000000000000000";
                  --when "000000000000000000000000000001" => output <= "00100100000000110000100000000000";
                  --when "000000000000000000000000000010" => output <= "00100100000001000001000000000000";
                  --when "000000000000000000000000000011" => output <= "10101100011000100000000000000000";
                  --when "000000000000000000000000000100" => output <= "00100000010000100000000000000001";
                  --when "000000000000000000000000000101" => output <= "00100000011000110000000000000100";
                  --when "000000000000000000000000000110" => output <= "00010100011001001111111111111100";
                  --when "000000000000000000000000000111" => output <= "00000000000000000000000000000000";
                  --when "000000000000000000000000001000" => output <= "00000000000000000000000000000000";
                  --when "000000000000000000000000001001" => output <= "00100100000000110000100000000000";
                  --when "000000000000000000000000001010" => output <= "10001100011000100000000000000000";
                  --when "000000000000000000000000001011" => output <= "00111100000000010000000000001000";
                  --when "000000000000000000000000001100" => output <= "10101100001000100000000000000000";
                  --when "000000000000000000000000001101" => output <= "00100000011000110000000000000100";
                  --when "000000000000000000000000001110" => output <= "00010100011001001111111111111011";
                  --when "000000000000000000000000001111" => output <= "00000000000000000000000000000000";
                  --when "000000000000000000000000010000" => output <= "00000000000000000000000000000000";
                  --when "000000000000000000000000010001" => output <= "00001000000000000000000000000000";
                  --when "000000000000000000000000010010" => output <= "00000000000000000000000000000000";
                  --when "000000000000000000000000010011" => output <= "00000000000000000000000000000000";

                  -- BOOT ROM - see boot.s
                  when "000000000000000000000000000000" => output <= "00111100000001000000000000001000";
                  when "000000000000000000000000000001" => output <= "10101100100000000000000000000000";
                  when "000000000000000000000000000010" => output <= "10101100100000000000000000000000";
                  when "000000000000000000000000000011" => output <= "10101100100000000000000000000000";
                  when "000000000000000000000000000100" => output <= "10101100100000000000000000000000";
                  when "000000000000000000000000000101" => output <= "00100100000000100000000001001101";
                  when "000000000000000000000000000110" => output <= "10101100100000100000000000000000";
                  when "000000000000000000000000000111" => output <= "00100100000000100000000001001001";
                  when "000000000000000000000000001000" => output <= "10101100100000100000000000000000";
                  when "000000000000000000000000001001" => output <= "00100100000000100000000001010000";
                  when "000000000000000000000000001010" => output <= "10101100100000100000000000000000";
                  when "000000000000000000000000001011" => output <= "00100100000000100000000001010011";
                  when "000000000000000000000000001100" => output <= "10101100100000100000000000000000";
                  when "000000000000000000000000001101" => output <= "00100100000000100000000000100000";
                  when "000000000000000000000000001110" => output <= "10101100100000100000000000000000";
                  when "000000000000000000000000001111" => output <= "00100100000000100000000001110010";
                  when "000000000000000000000000010000" => output <= "10101100100000100000000000000000";
                  when "000000000000000000000000010001" => output <= "00100100000000100000000001100101";
                  when "000000000000000000000000010010" => output <= "10101100100000100000000000000000";
                  when "000000000000000000000000010011" => output <= "00100100000000100000000001100001";
                  when "000000000000000000000000010100" => output <= "10101100100000100000000000000000";
                  when "000000000000000000000000010101" => output <= "00100100000000100000000001100100";
                  when "000000000000000000000000010110" => output <= "10101100100000100000000000000000";
                  when "000000000000000000000000010111" => output <= "00100100000000100000000001111001";
                  when "000000000000000000000000011000" => output <= "10101100100000100000000000000000";
                  when "000000000000000000000000011001" => output <= "00100100000000100000000000101110";
                  when "000000000000000000000000011010" => output <= "10101100100000100000000000000000";
                  when "000000000000000000000000011011" => output <= "00100000000000110000000000000000";
                  when "000000000000000000000000011100" => output <= "00111100000001111111111111111111";
                  when "000000000000000000000000011101" => output <= "00110100111001111111111111111111";
                  when "000000000000000000000000011110" => output <= "00100100000001010000000000000000";
                  when "000000000000000000000000011111" => output <= "10010000100001010000000000000100";
                  when "000000000000000000000000100000" => output <= "00000000000000000000000000000000";
                  when "000000000000000000000000100001" => output <= "00000000000001010010101000000000";
                  when "000000000000000000000000100010" => output <= "10010000100001100000000000000100";
                  when "000000000000000000000000100011" => output <= "00000000000000000000000000000000";
                  when "000000000000000000000000100100" => output <= "00000000101001100010100000100000";
                  when "000000000000000000000000100101" => output <= "00000000000001010010101000000000";
                  when "000000000000000000000000100110" => output <= "10010000100001100000000000000100";
                  when "000000000000000000000000100111" => output <= "00000000000000000000000000000000";
                  when "000000000000000000000000101000" => output <= "00000000101001100010100000100000";
                  when "000000000000000000000000101001" => output <= "00000000000001010010101000000000";
                  when "000000000000000000000000101010" => output <= "10010000100001100000000000000100";
                  when "000000000000000000000000101011" => output <= "00000000000000000000000000000000";
                  when "000000000000000000000000101100" => output <= "00000000101001100010100000100000";
                  when "000000000000000000000000101101" => output <= "10101100100000100000000000000000";
                  when "000000000000000000000000101110" => output <= "10101100011001010000000000000000";
                  when "000000000000000000000000101111" => output <= "00100000011000110000000000000100";
                  when "000000000000000000000000110000" => output <= "00010100101001111111111111101101";
                  when "000000000000000000000000110001" => output <= "00000000000000000000000000000000";
                  when "000000000000000000000000110010" => output <= "10101100011000001111111111111100";
                  when "000000000000000000000000110011" => output <= "10010000100001100000000000000100";
                  when "000000000000000000000000110100" => output <= "10010000100001100000000000000100";
                  when "000000000000000000000000110101" => output <= "10010000100001100000000000000100";
                  when "000000000000000000000000110110" => output <= "10010000100001100000000000000100";
                  when "000000000000000000000000110111" => output <= "10010000100001100000000000000100";
                  when "000000000000000000000000111000" => output <= "10010000100001100000000000000100";
                  when "000000000000000000000000111001" => output <= "10010000100001100000000000000100";
                  when "000000000000000000000000111010" => output <= "10010000100001100000000000000100";
                  when "000000000000000000000000111011" => output <= "00100100000000100000000001100111";
                  when "000000000000000000000000111100" => output <= "10101100100000100000000000000000";
                  when "000000000000000000000000111101" => output <= "00100100000000100000000001101111";
                  when "000000000000000000000000111110" => output <= "00001000000000000000000001000000";
                  when "000000000000000000000000111111" => output <= "10101100100000100000000000000000";

                  -- address not part of boot rom so give back sram content
                  when others => 
                     output <= sram_data_hi & sram_data_lo;
               end case;
	       
               -- recognize write cycle
               if mem_write = '1' then
		 mem_pause  <= '1';
		 next_state <= WRITE;
	       end if;

	       data <= sram_data_hi & sram_data_lo;

	    when WRITE =>
	       -- write correct data into memory
	       sram_we_hi <= mem_byte_sel(3) nor mem_byte_sel(2);
	       sram_we_lo <= mem_byte_sel(1) nor mem_byte_sel(0);

               if mem_byte_sel(3) = '1' then
	          sram_data_hi(15 downto 8) <= mem_data_w(31 downto 24);
	       else
	          sram_data_hi(15 downto 8) <= data(31 downto 24);
	       end if;

               if mem_byte_sel(2) = '1' then
                  sram_data_hi(7 downto 0) <= mem_data_w(23 downto 16);
               else
                  sram_data_hi(7 downto 0) <= data(23 downto 16);
               end if;

               if mem_byte_sel(1) = '1' then
                  sram_data_lo(15 downto 8) <= mem_data_w(15 downto 8);
               else
                  sram_data_lo(15 downto 8) <= data(15 downto 8);
               end if;

               if mem_byte_sel(0) = '1' then
                 sram_data_lo(7 downto 0) <= mem_data_w(7 downto 0);
               else
                  sram_data_lo(7 downto 0) <= data(7 downto 0);
               end if;

            when others => NULL;
	 end case;
      end if;
   end process; -- work

   mem_data_r   <= output;
end;


