---------------------------------------------------------------------
-- TITLE: Test Bench
-- AUTHOR: Steve Rhoads (rhoadss@yahoo.com)
-- DATE CREATED: 4/21/01
-- FILENAME: tbench.vhd
-- PROJECT: Plasma CPU core
-- COPYRIGHT: Software placed into the public domain by the author.
--    Software 'as is' without warranty.  Author liable for nothing.
-- DESCRIPTION:
--    This entity provides a test bench for testing the Plasma CPU core.
---------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use work.mlite_pack.all;

entity tbench is
end; --entity tbench

architecture logic of tbench is
   -- signals generated by testbench
   signal clk               : std_logic := '1';
   signal reset             : std_logic := '1';
   signal resetn            : std_logic;
   -- signals to uart
   signal TXD               : std_logic;
   signal RTS               : std_logic;
   signal CTS               : std_logic;
   signal CTS_ONE           : std_logic := '0';
   signal RXD               : std_logic;
   signal RXD_NULL          : std_logic := '1';
   -- signals to sram interface
   signal sram_we_hi        : std_logic;
   signal sram_we_lo        : std_logic;
   signal sram_ce_hi        : std_logic;
   signal sram_ce_lo        : std_logic;
   signal sram_oe_hi        : std_logic;
   signal sram_oe_lo        : std_logic;
   signal sram_address_hi   : std_logic_vector(18 downto 0);
   signal sram_address_lo   : std_logic_vector(18 downto 0);
   signal sram_data_hi      : std_logic_vector(15 downto 0);
   signal sram_data_lo      : std_logic_vector(15 downto 0);
   -- signals to mlite ram interface
   signal mem_byte_sel      : std_logic_vector(3 downto 0);
   signal mem_write         : std_logic;
   signal mem_address       : std_logic_vector(31 downto 0);
   signal mem_data_w        : std_logic_vector(31 downto 0);
   signal mem_data_r        : std_logic_vector(31 downto 0);
   -- signals to control second uart which outputs a test pattern
   signal uart_mem_byte_sel : std_logic_vector(3 downto 0) := "1111";
   signal uart_mem_write    : std_logic := '1';
   signal uart_mem_address  : std_logic_vector(31 downto 0) := "00000000000010000000000000000000";
   signal uart_mem_data_w   : std_logic_vector(31 downto 0) := "00000000000000000000000000100000";
   signal uart_mem_data_r   : std_logic_vector(31 downto 0);
   signal uart_mem_pause    : std_logic;
   signal uart_dbg          : std_logic_vector(7 downto 0);
begin  --architecture
   clk    <= not clk after 75 ns;
   reset  <= '0' after 1500 ns;
   resetn <= not reset;

   --Uncomment the line below to test interrupts
--   interrupt <= '1' after 20 us when interrupt = '0' else '0' after 400 ns;
   --Uncomment the line below to test mem_pause
--   mem_pause <= '1' after 100 ns when mem_pause = '0' else '0' after 100 ns;

   T1_cpu: plasma
      PORT MAP (
         BOARD_CLK       => clk,
         BOARD_RES       => resetn,

         BOARD_TXD       => TXD,
	 BOARD_RTS       => RTS,
	 BOARD_CTS       => CTS_ONE,
	 BOARD_RXD       => RXD_NULL,

         sram_we_hi      => sram_we_hi, 
         sram_we_lo      => sram_we_lo,
         sram_ce_hi      => sram_ce_hi,
         sram_ce_lo      => sram_ce_lo,
         sram_oe_hi      => sram_oe_hi,
         sram_oe_lo      => sram_oe_lo,
         sram_address_hi => sram_address_hi,
         sram_address_lo => sram_address_lo,
         sram_data_hi    => sram_data_hi,
         sram_data_lo    => sram_data_lo);

   T2_sram2mlite: sram2mlite
      PORT MAP (
         clk             => clk,

         mem_byte_sel    => mem_byte_sel,
         mem_write       => mem_write,
	 mem_address     => mem_address,
	 mem_data_w      => mem_data_w,
	 mem_data_r      => mem_data_r,

         sram_we_hi      => sram_we_hi,
         sram_we_lo      => sram_we_lo,
         sram_ce_hi      => sram_ce_hi,
         sram_ce_lo      => sram_ce_lo,
         sram_oe_hi      => sram_oe_hi,
         sram_oe_lo      => sram_oe_lo,
         sram_address_hi => sram_address_hi,
         sram_address_lo => sram_address_lo,
         sram_data_hi    => sram_data_hi,
         sram_data_lo    => sram_data_lo);

   T3_ram: ram
      PORT MAP (
         clk             => clk,
                                                                             
         mem_byte_sel    => mem_byte_sel,
         mem_write       => mem_write,
         mem_address     => mem_address,
         mem_data_w      => mem_data_w,
         mem_data_r      => mem_data_r);

   T4_uart: mlite2uart
      PORT MAP (
         reset           => reset,
	 clk             => clk,
	 mem_byte_sel    => uart_mem_byte_sel,
	 mem_write       => uart_mem_write,
	 mem_address     => uart_mem_address,
	 mem_data_w      => uart_mem_data_w,
	 mem_data_r      => uart_mem_data_r,
	 mem_pause       => uart_mem_pause,
	 TXD             => RXD,
	 RTS             => CTS,
	 CTS             => RTS,
	 RXD             => TXD,
	 dbg             => uart_dbg);

end; --architecture logic

