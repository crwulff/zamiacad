entity E5 is end; 

architecture arch of E5 is begin

end architecture;