entity top is
end entity top;


architecture RTL of top is
begin
  
  c0: entity WORK.COMP(RIGHTONE) ;
  
end architecture RTL;
