--------------------------------------------------------------------------
--  Crypto Chip
--  Copyright (C) 1999, Projektgruppe WS98/99
--  University of Stuttgart / Department of Computer Science / IFI-RA
--------------------------------------------------------------------------
-- Designer  : Thomas Stanka 
-- Group     : DES
--------------------------------------------------------------------
-- Design Unit Name : KEYVALID
-- Purpose : Part of the DES-module-core for the cryptochip "pg99"
-- 
-- File Name :  keyvalid.vhdl
--------------------------------------------------------------------
-- Simulator : SYNOPSYS VHDL System Simulator (VSS) Version 3.2.a
--------------------------------------------------------------------
-- Date 10.11.98   | Changes
--                 | 
--                 |
-----------------------------------------------------------------------

--------------------------------------------------------------------------
--  contents: this module checks for parity of an incomming key and creates 
--            secure keys when a key is created by random.
--------------------------------------------------------------------------
library IEEE;
   use IEEE.std_logic_1164.all;
   use IEEE.std_logic_arith.all; 

entity KEYVALID is
	port (KEY_IN : in  STD_LOGIC_VECTOR(63 downto 0);
	      KEY_OUT: out STD_LOGIC_VECTOR(55 downto 0);
              CTRL   : in  STD_LOGIC;                     -- has to be '0' if the key is generated by random
	      PARITY : out STD_LOGIC                      -- PARITY='1' <=> key has a false parity
	     );
end KEYVALID;

architecture BEHAVIORAL of KEYVALID is
begin
  process(KEY_IN,CTRL)
        variable PARITY_CHECK:STD_LOGIC_VECTOR(7 downto 0);
	begin	 

          -- first check the incoming key parity and send a warning over the parity-bit

	  PARITY_CHECK(0):= KEY_IN(0) xor KEY_IN(1) xor KEY_IN(2) xor KEY_IN(3) xor KEY_IN(4) xor KEY_IN(5) xor KEY_IN(6);
	  PARITY_CHECK(1):= KEY_IN(8) xor KEY_IN(9) xor KEY_IN(10) xor KEY_IN(11) xor KEY_IN(12) xor KEY_IN(13) xor KEY_IN(14);
	  PARITY_CHECK(2):= KEY_IN(16) xor KEY_IN(17) xor KEY_IN(18) xor KEY_IN(19) xor KEY_IN(20) xor KEY_IN(21) xor KEY_IN(22);
      	  PARITY_CHECK(3):= KEY_IN(24) xor KEY_IN(25) xor KEY_IN(26) xor KEY_IN(27) xor KEY_IN(28) xor KEY_IN(29) xor KEY_IN(30);
      	  PARITY_CHECK(4):= KEY_IN(32) xor KEY_IN(33) xor KEY_IN(34) xor KEY_IN(35) xor KEY_IN(36) xor KEY_IN(37) xor KEY_IN(38);
      	  PARITY_CHECK(5):= KEY_IN(40) xor KEY_IN(41) xor KEY_IN(42) xor KEY_IN(43) xor KEY_IN(44) xor KEY_IN(45) xor KEY_IN(46);
      	  PARITY_CHECK(6):= KEY_IN(48) xor KEY_IN(49) xor KEY_IN(50) xor KEY_IN(51) xor KEY_IN(52) xor KEY_IN(53) xor KEY_IN(54);
      	  PARITY_CHECK(7):= KEY_IN(56) xor KEY_IN(57) xor KEY_IN(58) xor KEY_IN(59) xor KEY_IN(60) xor KEY_IN(61) xor KEY_IN(62);
          parity<=(PARITY_CHECK(0) xor KEY_IN(7)) or (PARITY_CHECK(1) xor KEY_IN(15)) or (PARITY_CHECK(2) xor KEY_IN(23)) 
	       or (PARITY_CHECK(3) xor KEY_IN(31)) or (PARITY_CHECK(4) xor KEY_IN(39)) or (PARITY_CHECK(5) xor KEY_IN(47))
	       or (PARITY_CHECK(6) xor KEY_IN(55)) or (PARITY_CHECK(7) xor KEY_IN(63));   
	  
	  KEY_OUT( 6 downto  0) <= KEY_IN( 7 downto  1);
          KEY_OUT(13 downto  7) <= KEY_IN(15 downto  9);
          KEY_OUT(20 downto 14) <= KEY_IN(23 downto 17);
          KEY_OUT(27 downto 21) <= KEY_IN(31 downto 25);
          KEY_OUT(34 downto 28) <= KEY_IN(39 downto 33);
          KEY_OUT(41 downto 35) <= KEY_IN(47 downto 41);
          KEY_OUT(48 downto 42) <= KEY_IN(55 downto 49);
          KEY_OUT(55 downto 49) <= KEY_IN(63 downto 57);  
          
          -- if the key is generated by random then set bit 1 and 2 to "01" in order to get secure keys
	  -- this reduces the keyspace to 25% but it's safty and fast to go
 	  if CTRL='0' then
          	  KEY_OUT(1 downto 0)<="10";
	  end if; 

	end process;

end BEHAVIORAL;



