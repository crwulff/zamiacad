-------------------------------------------------------------------------------
-- Title      : Initialized On Chip Sync RAM
-- Description: Auto Created by gen_vhdl_ram from manikremote.bin
-------------------------------------------------------------------------------
-- File       : manikremote.vhd
-- Author     : gen_vhdl_mem
-- Company    : NikTech Inc.
-- Created    : Mon Oct  9 21:26:38 2006

-------------------------------------------------------------------------------
-- Copyright (c) 2005 
-------------------------------------------------------------------------------
-------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
entity manikremote is
generic (WIDTH      : integer := 32;
         ADDR_WIDTH : integer := 32);
port (clk   : std_logic;
reset : std_logic;
-- Wishbone slave interface
WBS_ADR_I : in  std_logic_vector (ADDR_WIDTH-1 downto 0);
WBS_SEL_I : in  std_logic_vector (3 downto 0);
WBS_DAT_I : in  std_logic_vector (WIDTH-1 downto 0);
WBS_WE_I  : in  std_logic;
WBS_STB_I : in  std_logic;
WBS_CYC_I : in  std_logic;
WBS_CTI_I : in  std_logic_vector (2 downto 0);
WBS_BTE_I : in  std_logic_vector (1 downto 0);
WBS_DAT_O : out std_logic_vector (WIDTH-1 downto 0);
WBS_ACK_O : out std_logic;
WBS_ERR_O : out std_logic);
end manikremote;
architecture RTL of manikremote is
signal ben : std_logic_vector (3 downto 0) := "0000";
signal wen : std_logic_vector (3 downto 0) := "0000";
signal ack : std_logic := '0';
begin
ben(0) <= WBS_STB_I and WBS_SEL_I(3);
ben(1) <= WBS_STB_I and WBS_SEL_I(2);
ben(2) <= WBS_STB_I and WBS_SEL_I(1);
ben(3) <= WBS_STB_I and WBS_SEL_I(0);
wen(0) <= WBS_WE_I and WBS_STB_I and WBS_SEL_I(3);
wen(1) <= WBS_WE_I and WBS_STB_I and WBS_SEL_I(2);
wen(2) <= WBS_WE_I and WBS_STB_I and WBS_SEL_I(1);
wen(3) <= WBS_WE_I and WBS_STB_I and WBS_SEL_I(0);
process (clk, reset)
begin
if reset = '1' then
ack <= '0';
elsif rising_edge(clk) then
if ack = '1' then
ack <= '0' after 1 ns;
else
ack <= WBS_STB_I after 1 ns;
end if;
end if;
end process;
WBS_ACK_O <= ack;
WBS_ERR_O <= '0';
mem_block: block
signal raddr,waddr : std_logic_vector (8-1 downto 0) := (others => '0');
signal data_int    : std_logic_vector (WIDTH-1 downto 0);
signal data_w      : std_logic_vector (WIDTH-1 downto 0);
signal we          : std_logic := '0' ;
type ram_mem_type is array(0 to 256-1) of std_logic_vector(32-1 downto 0);
attribute syn_ramstyle : string;
signal ram_mem0 : ram_mem_type := (
"11110000000000000000000000001001", -- 0xf0000009 0x0
"11110000000000000000000001000110", -- 0xf0000046 0x4
"11110000000000000000000000101100", -- 0xf000002c 0x8
"11110000000000000000000000110110", -- 0xf0000036 0xc
"11110000000000000000000000000101", -- 0xf0000005 0x10
"01000011000010010111000000010000", -- 0x43097010 0x14
"00010011000000010001000000001111", -- 0x1301100f 0x18
"11110100001110110001001011110010", -- 0xf43b12f2 0x1c
"10010001111100000001001011110010", -- 0x91f012f2 0x20
"10010100111100000001001011110011", -- 0x94f012f3 0x24
"10010101111100000001001011110110", -- 0x95f012f6 0x28
"10010110111100000001001011110111", -- 0x96f012f7 0x2c
"10010111111100000001001011111000", -- 0x97f012f8 0x30
"10011000111100000001001011111001", -- 0x98f012f9 0x34
"10011001111100000001001011111010", -- 0x99f012fa 0x38
"10011010111100001000000011110000", -- 0x9af080f0 0x3c
"01101100000001001001000000000000", -- 0x6c049000 0x40
"10010001000100001001001000100000", -- 0x91109220 0x44
"10010011001100001001010001000000", -- 0x93309440 0x48
"10010101010100001001011001100000", -- 0x95509660 0x4c
"10010111011100001001100010000000", -- 0x97709880 0x50
"10011001100100001001101010100000", -- 0x99909aa0 0x54
"10011011101100001001110011000000", -- 0x9bb09cc0 0x58
"10011101110100001001111011100000", -- 0x9dd09ee0 0x5c
"00011110000000010110110100000100", -- 0x1e016d04 0x60
"10010000111100000001001011110000", -- 0x90f012f0 0x64
"10010010111100000001001011110001", -- 0x92f012f1 0x68
"10010011111100001111101111111111", -- 0x93f0fbff 0x6c
"11111111110101110010010000010000", -- 0xffd72410 0x70
"11111000000000000000000001000101", -- 0xf8000045 0x74
"11110100000110110110110100000100", -- 0xf41b6d04 0x78
"10010000111100000001001011110000", -- 0x90f012f0 0x7c
"10010010111100000001001011110001", -- 0x92f012f1 0x80
"10010011111100001111101111111111", -- 0x93f0fbff 0x84
"11111111110010110010010000010000", -- 0xffcb2410 0x88
"11111000000000000000000100101001", -- 0xf8000129 0x8c
"11110100000011110110110100000100", -- 0xf40f6d04 0x90
"10010000111100000001001011110000", -- 0x90f012f0 0x94
"10010010111100000001001011110001", -- 0x92f012f1 0x98
"10010011111100001111101111111111", -- 0x93f0fbff 0x9c
"11111111101111110010011100010001", -- 0xffbf2711 0xa0
"00010011011000010010010000010000", -- 0x13612410 0xa4
"11111000000000000000000010000011", -- 0xf8000083 0xa8
"11110100000000011000000100010000", -- 0xf4018110 0xac
"10000010001000001000001100110000", -- 0x82208330 0xb0
"10000100010000001000010101010000", -- 0x84408550 0xb4
"10000110011000001000011101110000", -- 0x86608770 0xb8
"10001000100000001000100110010000", -- 0x88808990 0xbc
"10001010101000001000101110110000", -- 0x8aa08bb0 0xc0
"10001100110000001000110111010000", -- 0x8cc08dd0 0xc4
"10001110111000000110001100001100", -- 0x8ee0630c 0xc8
"10001010111100000001001110101111", -- 0x8af013af 0xcc
"10001001111100000001001110011111", -- 0x89f0139f 0xd0
"10001000111100000001001110001111", -- 0x88f0138f 0xd4
"10000111111100000001001101111111", -- 0x87f0137f 0xd8
"10000110111100000001001101101111", -- 0x86f0136f 0xdc
"10000100111100000001001100101111", -- 0x84f0132f 0xe0
"10000011111100000001001100011111", -- 0x83f0131f 0xe4
"10000010111100000001001100001111", -- 0x82f0130f 0xe8
"10000001111100000001001100101111", -- 0x81f0132f 0xec
"10000000111100000110001000001100", -- 0x80f0620c 0xf0
"00011110000000100000000000000000", -- 0x1e020000 0xf4
"00000000000000000000001111111000", -- 0x000003f8 0xf8
"00100100000000000010010000000000", -- 0x24002400 0xfc
"01101111000011000001001001010001", -- 0x6f0c1251 0x100
"10010000010100000100000001110100", -- 0x90504074 0x104
"10000000011101110011000001110000", -- 0x80773070 0x108
"11101100000000110001110100000111", -- 0xec031d07 0x10c
"00000000000000001000000001010000", -- 0x00008050 0x110
"01100000000001000001110000000101", -- 0x60041c05 0x114
"00000000000000000000001101011100", -- 0x0000035c 0x118
"00100100000000000010010000000000", -- 0x24002400 0x11c
"01101111000001000001001001010001", -- 0x6f041251 0x120
"10010000111100001001000111100000", -- 0x90f091e0 0x124
"10010010010100000010010011100010", -- 0x925024e2 0x128
"00100100111100010110111111111111", -- 0x24f16fff 0x12c
"00110000111111111110110000001110", -- 0x30ffec0e 0x130
"00010010011100000100000001101000", -- 0x12704068 0x134
"00100110011101100001001100000111", -- 0x26761307 0x138
"11000000000111101111100000000000", -- 0xc01ef800 0x13c
"00000001000000000110000011100001", -- 0x010060e1 0x140
"00010010011100000100000001100101", -- 0x12704065 0x144
"00100101011101100001001100000111", -- 0x25761307 0x148
"11110111111100011000000011110000", -- 0xf7f180f0 0x14c
"10000001111000001000001001010000", -- 0x81e08250 0x150
"01100000000011000001110000000101", -- 0x600c1c05 0x154
"00000000000000000000010000000000", -- 0x00000400 0x158
"11111111111111111111101111111111", -- 0xfffffbff 0x15c
"01101111000001001001000011110000", -- 0x6f0490f0 0x160
"00010010010100011001000111100000", -- 0x125191e0 0x164
"00100100111100011001001001010000", -- 0x24f19250 0x168
"00100100111000100111010000011101", -- 0x24e2741d 0x16c
"11111000000000000000000011100111", -- 0xf80000e7 0x170
"01101111111111110011000011111111", -- 0x6fff30ff 0x174
"11101100000011111111100000000000", -- 0xec0ff800 0x178
"00000000111010100101111100011111", -- 0x00ea5f1f 0x17c
"00010010011100000100000001100111", -- 0x12704067 0x180
"00100110011101100001001100000111", -- 0x26761307 0x184
"11010000000111100110000011100001", -- 0xd01e60e1 0x188
"00010010011100000100000001100101", -- 0x12704065 0x18c
"00100101011101100001001100000111", -- 0x25761307 0x190
"11110111111100001000000011110000", -- 0xf7f080f0 0x194
"10000001111000001000001001010000", -- 0x81e08250 0x198
"01100000000011000001110000000101", -- 0x600c1c05 0x19c
"00000000000000000000100000000000", -- 0x00000800 0x1a0
"11111111111111111111011111111111", -- 0xfffff7ff 0x1a4
"00100100000000000010010000000000", -- 0x24002400 0x1a8
"00100100000000000010010000000000", -- 0x24002400 0x1ac
"01101110000001001001010010110000", -- 0x6e0494b0 0x1b0
"10010011110000000001001001010001", -- 0x93c01251 0x1b4
"00100100101100011001010110100000", -- 0x24b195a0 0x1b8
"10010000111100001001000111100000", -- 0x90f091e0 0x1bc
"10010010110100001001011001010000", -- 0x92d09650 0x1c0
"00100100110000010110010010110100", -- 0x24c164b4 0x1c4
"10000000111110110111000000010001", -- 0x80fb7011 0x1c8
"11111000000000000000000010110001", -- 0xf80000b1 0x1cc
"00100100011111110101000001110001", -- 0x247f5071 0x1d0
"01110000101000000011000001110000", -- 0x70a03070 0x1d4
"11101100000101110010100101111111", -- 0xec17297f 0x1d8
"00101011011101110101000001111111", -- 0x2b77507f 0x1dc
"00110000011100011110010000010010", -- 0x3071e412 0x1e0
"10000001011111000011000001110010", -- 0x817c3072 0x1e4
"11100100000000110100001101111010", -- 0xe403437a 0x1e8
"11110100000010000011000001110011", -- 0xf4083073 0x1ec
"11100100011000101000001101111100", -- 0xe462837c 0x1f0
"00100001011101110010000101110111", -- 0x21772177 0x1f4
"01000011011010000010000101110110", -- 0x43682176 0x1f8
"10000000010101111000001001101100", -- 0x8057826c 0x1fc
"10010000011001111001000101011100", -- 0x9067915c 0x200
"11110100010110000111010100011000", -- 0xf4587518 0x204
"11111000000000000000000010011011", -- 0xf800009b 0x208
"11111000000000000000000010100001", -- 0xf80000a1 0x20c
"00100100111000010101111111101111", -- 0x24e15fef 0x210
"01110110011100110011000111100111", -- 0x767331e7 0x214
"11101100010010000111011001110100", -- 0xec487674 0x218
"00110100111001111110010000000110", -- 0x34e7e406 0x21c
"01110100011111010011000111100111", -- 0x747d31e7 0x220
"11101100000010100111010101110010", -- 0xec0a7572 0x224
"11110100000001010111011001111101", -- 0xf405767d 0x228
"00110001111001111110110000000101", -- 0x31e7ec05 0x22c
"01110111011100100011000111100111", -- 0x777231e7 0x230
"11101100001001101111010000111010", -- 0xec26f43a 0x234
"11111000000000000000000010001011", -- 0xf800008b 0x238
"00100100110100011111100000000000", -- 0x24d1f800 0x23c
"00000000100010000101111111011111", -- 0x00885fdf 0x240
"01011111000111110000110011011000", -- 0x5f1f0cd8 0x244
"00100110110100011111100000000000", -- 0x26d1f800 0x248
"00000000100000100010010011110001", -- 0x008224f1 0x24c
"11111000000000000000000001111111", -- 0xf800007f 0x250
"01011111111111110101111100011111", -- 0x5fff5f1f 0x254
"00001100111110000010011011110001", -- 0x0cf826f1 0x258
"11111000000000000000000001111001", -- 0xf8000079 0x25c
"01011111000111110000110011111000", -- 0x5f1f0cf8 0x260
"00100110111100011111100000000000", -- 0x26f1f800 0x264
"00000000011101000000110011111000", -- 0x00740cf8 0x268
"01011111000111110111011001111101", -- 0x5f1f767d 0x26c
"00100110111100010011000111100111", -- 0x26f131e7 0x270
"00111100000111010011110000101111", -- 0x3c1d3c2f 0x274
"11101100000011110010010000011101", -- 0xec0f241d 0x278
"00100100001011111111010000010010", -- 0x242ff412 0x27c
"11111000000000000000000001100111", -- 0xf8000067 0x280
"01011111000111110111011101110010", -- 0x5f1f7772 0x284
"00110001111001110010000100010001", -- 0x31e72111 0x288
"00100001000100011110010000000111", -- 0x2111e407 0x28c
"00100100001011000010000100100001", -- 0x242c2121 0x290
"01110000000101001111101111111111", -- 0x7014fbff 0x294
"11111111010001001111010000001000", -- 0xff44f408 0x298
"00100100001011000010000100100001", -- 0x242c2121 0x29c
"01110000000101001111101111111111", -- 0x7014fbff 0x2a0
"11111111010111101111010000000010", -- 0xff5ef402 0x2a4
"01110000101000010111011000011011", -- 0x70a1761b 0x2a8
"11111000000000000000000001001001", -- 0xf8000049 0x2ac
"00110000101000001110111110101101", -- 0x30a0efad 0x2b0
"10000000011110110100000001101001", -- 0x807b4069 0x2b4
"00100110011101101001000001111011", -- 0x2676907b 0x2b8
"10000110010100001000000011110000", -- 0x865080f0 0x2bc
"10000001111000001000001011010000", -- 0x81e082d0 0x2c0
"10000011110000001000010010110000", -- 0x83c084b0 0x2c4
"10000101101000000111000000010000", -- 0x85a07010 0x2c8
"00010011000101010110000100001100", -- 0x1315610c 0x2cc
"11110000000000000000000000101111", -- 0xf000002f 0x2d0
"00000000000000000000001101011100", -- 0x0000035c 0x2d4
"00000000000000000000001101100000", -- 0x00000360 0x2d8
"00000000000100000000000000100000", -- 0x00100020 0x2dc
"01101111000011000001001001010001", -- 0x6f0c1251 0x2e0
"10010000010100000100000100110000", -- 0x90504130 0x2e4
"01110000010000000010010001010100", -- 0x70402454 0x2e8
"01000001011100000010010001100001", -- 0x41702461 0x2ec
"00100001010101010010000101010101", -- 0x21552155 0x2f0
"01100100011001000010000101010111", -- 0x64642157 0x2f4
"10000000011101100010010101110011", -- 0x80762573 0x2f8
"00100001001100110011000001110000", -- 0x21333070 0x2fc
"11101100000011100011000001000000", -- 0xec0e3040 0x300
"11100100000001101000000001010000", -- 0xe4068050 0x304
"00010011000101010110000000000100", -- 0x13156004 0x308
"11110011111111111111111101010001", -- 0xf3ffff51 0x30c
"10000000011101010011000001110000", -- 0x80753070 0x310
"11101100000001000001110100000111", -- 0xec041d07 0x314
"00000000000000001111010000000100", -- 0x0000f404 0x318
"01100000010000010011011001000110", -- 0x60413646 0x31c
"11101111111001011000000001010000", -- 0xefe58050 0x320
"01100000000001000001110000000101", -- 0x60041c05 0x324
"00000100000000000000000000000000", -- 0x04000000 0x328
"00000000000000000000001101100000", -- 0x00000360 0x32c
"00110000000100001110110000000010", -- 0x3010ec02 0x330
"01110001000100000100000001110001", -- 0x71104071 0x334
"11010000000101110001111000000001", -- 0xd0171e01 0x338
"10000000000000000000000000000001", -- 0x80000001 0x33c
"01000000011100101101000000010111", -- 0x4072d017 0x340
"00011110000000010000000000000000", -- 0x1e010000 0x344
"10000000000000000000000000000000", -- 0x80000000 0x348
"00100100000000000010010000000000", -- 0x24002400 0x34c
"01000000000100101100000000010001", -- 0x4012c011 0x350
"00011110000000010000000000000000", -- 0x1e010000 0x354
"10000000000000000000000000000000", -- 0x80000000 0x358
"00000000000000000000000000000000", -- 0x00000000 0x35c
"00000000000000000000000000000000", -- 0x00000000 0x360
"00000000000000000000000000000000", -- 0x00000000 0x364
"00000000000000000000000000000000", -- 0x00000000 0x368
"00000000000000000000000000000000", -- 0x00000000 0x36c
"00000000000000000000000000000000", -- 0x00000000 0x370
"00000000000000000000000000000000", -- 0x00000000 0x374
"00000000000000000000000000000001", -- 0x00000001 0x378
"00000000000000000000000000000000", -- 0x00000000 0x37c
"00000000000000000000000000000000", -- 0x00000000 0x380
"00000000000000000000000000000000", -- 0x00000000 0x384
"00000000000000000000000000000000", -- 0x00000000 0x388
"00000000000000000000000000000000", -- 0x00000000 0x38c
"00000000000000000000000000000000", -- 0x00000000 0x390
"00000000000000000000000000000000", -- 0x00000000 0x394
"00000000000000000000000000000000", -- 0x00000000 0x398
"00000000000000000000000000000000", -- 0x00000000 0x39c
"00000000000000000000000000000000", -- 0x00000000 0x3a0
"00000000000000000000000000000000", -- 0x00000000 0x3a4
"00000000000000000000000000000000", -- 0x00000000 0x3a8
"00000000000000000000000000000000", -- 0x00000000 0x3ac
"00000000000000000000000000000000", -- 0x00000000 0x3b0
"00000000000000000000000000000000", -- 0x00000000 0x3b4
"00000000000000000000000000000000", -- 0x00000000 0x3b8
"00000000000000000000000000000000", -- 0x00000000 0x3bc
"00000000000000000000000000000000", -- 0x00000000 0x3c0
"00000000000000000000000000000000", -- 0x00000000 0x3c4
"00000000000000000000000000000000", -- 0x00000000 0x3c8
"00000000000000000000000000000000", -- 0x00000000 0x3cc
"00000000000000000000000000000000", -- 0x00000000 0x3d0
"00000000000000000000000000000000", -- 0x00000000 0x3d4
"00000000000000000000000000000000", -- 0x00000000 0x3d8
"00000000000000000000000000000000", -- 0x00000000 0x3dc
"00000000000000000000000000000000", -- 0x00000000 0x3e0
"00000000000000000000000000000000", -- 0x00000000 0x3e4
"00000000000000000000000000000000", -- 0x00000000 0x3e8
"00000000000000000000000000000000", -- 0x00000000 0x3ec
"00000000000000000000000000000000", -- 0x00000000 0x3f0
"00000000000000000000000000000000", -- 0x00000000 0x3f4
"00000000000000000000000000000000", -- 0x3f8
"00000000000000000000000000000000" -- 0x3fc
);
attribute syn_ramstyle of ram_mem0 : signal is "block_ram";
begin
process (clk)
begin
if rising_edge(clk) then
raddr <= WBS_ADR_I(8+1 downto 2);
end if;
end process;
waddr <= WBS_ADR_I(8+1 downto 2);
process (clk, reset)
begin
if reset = '1' then
we    <= '0';
elsif rising_edge(clk) then
if WBS_STB_I = '1' and WBS_WE_I = '1'  and ack = '0' then
we <= '1';
else
we <= '0';
end if;
end if;
end process ;
process (clk)
begin
if rising_edge(clk) then
if we = '1' then
ram_mem0(conv_integer(waddr)) <= data_w((WIDTH*1/1)-1 downto WIDTH*0/1);
end if;
end if;
end process ;
data_int <= ram_mem0(conv_integer(raddr));
data_w(WIDTH-1 downto 3*WIDTH/4) <= WBS_DAT_I(WIDTH-1 downto 3*WIDTH/4) when WBS_SEL_I(3) = '1' else
data_int(WIDTH-1 downto 3*WIDTH/4); 
data_w((3*WIDTH/4)-1 downto 2*WIDTH/4) <= WBS_DAT_I((3*WIDTH/4)-1 downto 2*WIDTH/4) when WBS_SEL_I(2)='1' else
data_int((3*WIDTH/4)-1 downto 2*WIDTH/4); 
data_w((2*WIDTH/4)-1 downto 1*WIDTH/4) <= WBS_DAT_I((2*WIDTH/4)-1 downto 1*WIDTH/4) when WBS_SEL_I(1)='1' else
data_int((2*WIDTH/4)-1 downto 1*WIDTH/4); 
data_w((1*WIDTH/4)-1 downto 0*WIDTH/4) <= WBS_DAT_I((1*WIDTH/4)-1 downto 0*WIDTH/4) when WBS_SEL_I(0)='1' else
data_int((1*WIDTH/4)-1 downto 0*WIDTH/4); 
WBS_DAT_O <= data_int;
end block mem_block ;
end RTL;
