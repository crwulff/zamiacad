-- VHDL Model Created from SGE Symbol fsm.sym -- Jan  4 19:36:28 1999

--------------------------------------------------------------------------
----------------------------------------------------------------------
--  Crypto Chip
--  Copyright (C) 1999, Projektgruppe WS98/99
--  University of Stuttgart / Department of Computer Science / IFI-RA
--------------------------------------------------------------------------
-- Designers : Jens Kuenzer
-- Group     : CTRL
--------------------------------------------------------------------
-- Design Unit Name : FSM
-- Purpose : Steuerwerk fuer das main_ctrl
-- 
-- File Name : fsm.vhd
--------------------------------------------------------------------
-- Simulator : SYNOPSYS VHDL System Simulator (VSS) Version 3.2.a
--------------------------------------------------------------------
-- Date  24.11.98  | Changes
--       09.12.98  | begin with debug
--       14.12.98  | RSA tested with success
--	 15.12.98  | read-data&keys functionality added
--       04.01.98  | check authentify testable
--		   | ENABLE_TEST pin added
-----------------------------------------------------------------------

--------------------------------------------------------------------------
--  Ein grosser endlicher Automat um alles zu steuern.
--  und ein 8 Bit Zaehler
--------------------------------------------------------------------------
library IEEE;
   use IEEE.std_logic_1164.all;
   use IEEE.std_logic_misc.all;
package RAM_ADR_CONST is
    constant RSAKEYSIZE		: STD_LOGIC_VECTOR(7 downto 0) := "00011000";
    constant RAM_ADR_PUBLICKEY	: STD_LOGIC_VECTOR(7 downto 0) := "00000000";
    constant RAM_ADR_PRIVATKEY	: STD_LOGIC_VECTOR(7 downto 0) := "00011000";
    constant RAM_ADR_MODUL	: STD_LOGIC_VECTOR(7 downto 0) := "00110000";
    constant RAM_ADR_ZERT	: STD_LOGIC_VECTOR(7 downto 0) := "01001000";
    constant RAM_ADR_ZERTPUB	: STD_LOGIC_VECTOR(7 downto 0) := "01100000";
    constant RAM_ADR_ZERTMODUL	: STD_LOGIC_VECTOR(7 downto 0) := "01111000";
    constant RAM_ADR_TEMPEXP    : STD_LOGIC_VECTOR(7 downto 0) := "10010000";
    constant RAM_ADR_PIN	: STD_LOGIC_VECTOR(7 downto 0) := "10101000";
    constant RAM_ADR_DES_KEY	: STD_LOGIC_VECTOR(7 downto 0) := "10101001";
    constant RAM_ADR_USER	: STD_LOGIC_VECTOR(7 downto 0) := "10101011";

    constant RAM_MODE_NOP		: STD_LOGIC_VECTOR(5 downto 0) := "000000";
    constant RAM_MODE_INC		: STD_LOGIC_VECTOR(5 downto 0) := "100000";
    constant RAM_MODE_SET_PUBLICKEY	: STD_LOGIC_VECTOR(5 downto 0) := "010000";
    constant RAM_MODE_SET_PRIVATKEY	: STD_LOGIC_VECTOR(5 downto 0) := "010110";
    constant RAM_MODE_SET_MODUL		: STD_LOGIC_VECTOR(5 downto 0) := "010001";
    constant RAM_MODE_SET_ZERT		: STD_LOGIC_VECTOR(5 downto 0) := "010100";
    constant RAM_MODE_SET_ZERTPUB	: STD_LOGIC_VECTOR(5 downto 0) := "010111";
    constant RAM_MODE_SET_ZERTMODUL	: STD_LOGIC_VECTOR(5 downto 0) := "010010";
    constant RAM_MODE_SET_TEMPEXP	: STD_LOGIC_VECTOR(5 downto 0) := "011110";
    constant RAM_MODE_SET_PIN		: STD_LOGIC_VECTOR(5 downto 0) := "011100";
    constant RAM_MODE_SET_DES_KEY	: STD_LOGIC_VECTOR(5 downto 0) := "011101";
    constant RAM_MODE_SET_USER		: STD_LOGIC_VECTOR(5 downto 0) := "011111";
end RAM_ADR_CONST;

library IEEE;
   use IEEE.std_logic_1164.all;
   use IEEE.std_logic_misc.all;
   use IEEE.std_logic_arith.all;
   use IEEE.std_logic_unsigned.all;
   use WORK.RAM_ADR_CONST.all;

-- purpose: Calculates(set and count) the RAM-adress.
entity RAM_COUNTER is
    port ( RAM_ADR : out STD_LOGIC_VECTOR(7 downto 0);
	   CLK : in STD_LOGIC;  	-- clock
	   RESET : in STD_LOGIC;  	-- reset
	   RAM_MODE : in STD_LOGIC_VECTOR(5 downto 0);
	   RAM_ADR_IS_AT_END_OFF_ALL		: Out   std_logic;
	   RAM_ADR_IS_AT_END_OFF_TEMPEXP	: Out   std_logic;
	   RAM_ADR_IS_AT_END_OFF_MODUL		: Out   std_logic;
	   RAM_ADR_IS_AT_END_OFF_PUBLICKEY	: Out   std_logic;
	   RAM_ADR_IS_AT_END_OFF_PRIVATKEY	: Out   std_logic;
	   RAM_ADR_IS_AT_END_OFF_ZERTPUB	: Out   std_logic;
	   RAM_ADR_IS_AT_END_OFF_ZERTMODUL	: Out   std_logic;
	   INVERT : in STD_LOGIC );
end RAM_COUNTER;

architecture BEHAVIORAL of RAM_COUNTER is
    
    signal RAM_ADR_I : STD_LOGIC_VECTOR(7 downto 0);
    
begin  -- RAM_COUNTER

    -- purpose: Calculates(set and count) the RAM-adress.
    -- type:    memorizing
    -- inputs:  CLK, RESET, RAM_MODE, RAM_ADR_I
    -- outputs: RAM_ADR_I
    P_RAM_ADR : process (CLK, RESET)
    begin
	-- activities triggered by asynchronous reset (active high)
	if RESET = '1' then
	    RAM_ADR_I <= (others => '0');
	-- activities triggered by rising edge of clock
	elsif CLK'event and CLK = '1' then
	    case RAM_MODE is
		when RAM_MODE_INC =>
		    RAM_ADR_I <= RAM_ADR_I + "00000001";
		when RAM_MODE_SET_PRIVATKEY =>
		    RAM_ADR_I <= RAM_ADR_PRIVATKEY;
		when RAM_MODE_SET_PUBLICKEY =>
		    RAM_ADR_I <= RAM_ADR_PUBLICKEY;
		when RAM_MODE_SET_TEMPEXP =>
		    RAM_ADR_I <= RAM_ADR_TEMPEXP;
		when RAM_MODE_SET_ZERTMODUL =>
		    RAM_ADR_I <= RAM_ADR_ZERTMODUL;
		when RAM_MODE_SET_ZERTPUB =>
		    RAM_ADR_I <= RAM_ADR_ZERTPUB;
		when RAM_MODE_SET_ZERT =>
		    RAM_ADR_I <= RAM_ADR_ZERT;
		when RAM_MODE_SET_USER =>
		    RAM_ADR_I <= RAM_ADR_USER;
		when RAM_MODE_SET_DES_KEY =>
		    RAM_ADR_I <= RAM_ADR_DES_KEY;
		when RAM_MODE_SET_MODUL =>
		    RAM_ADR_I <= RAM_ADR_MODUL;
		when RAM_MODE_SET_PIN =>
		    RAM_ADR_I <= RAM_ADR_PIN;
		when others => NULL;
	    end case;
	end if;
    end process P_RAM_ADR;

    RAM_ADR <= not RAM_ADR_I when INVERT = '1' else RAM_ADR_I;

    process (RAM_ADR_I)	
    begin  -- process
	   RAM_ADR_IS_AT_END_OFF_ALL <= '0'; 
	   RAM_ADR_IS_AT_END_OFF_TEMPEXP <= '0'; 
	   RAM_ADR_IS_AT_END_OFF_MODUL <= '0'; 
	   RAM_ADR_IS_AT_END_OFF_PUBLICKEY <= '0'; 
	   RAM_ADR_IS_AT_END_OFF_PRIVATKEY <= '0'; 
	   RAM_ADR_IS_AT_END_OFF_ZERTPUB <= '0'; 
	   RAM_ADR_IS_AT_END_OFF_ZERTMODUL <= '0';
	
	if RAM_ADR_I = RAM_ADR_PUBLICKEY then
	   RAM_ADR_IS_AT_END_OFF_ALL <= '1'; 
	end if;
	if RAM_ADR_I = RAM_ADR_PIN then
	   RAM_ADR_IS_AT_END_OFF_TEMPEXP <= '1'; 
	end if;
	if RAM_ADR_I = RAM_ADR_ZERT then
	   RAM_ADR_IS_AT_END_OFF_MODUL <= '1'; 
	end if;
	if RAM_ADR_I = RAM_ADR_PRIVATKEY then
	   RAM_ADR_IS_AT_END_OFF_PUBLICKEY <= '1'; 
	end if;
	if RAM_ADR_I = RAM_ADR_MODUL then
	   RAM_ADR_IS_AT_END_OFF_PRIVATKEY <= '1'; 
	end if;
	if RAM_ADR_I = RAM_ADR_ZERTMODUL then
	   RAM_ADR_IS_AT_END_OFF_ZERTPUB <= '1'; 
	end if;
	if RAM_ADR_I = RAM_ADR_TEMPEXP then
	   RAM_ADR_IS_AT_END_OFF_ZERTMODUL <= '1';
	end if;
    end process;
    
end BEHAVIORAL;


library IEEE;
   use IEEE.std_logic_1164.all;
   use IEEE.std_logic_misc.all;
   use WORK.RAM_ADR_CONST.all;

entity FSM_CORE is
      Port ( CARDCHANGE : In    std_logic;
	     CLK : In    std_logic;
	     CTRL : In    std_logic_vector (7 downto 0);
             CTRL_CHANGE : In    std_logic;
             DATA_VALID : In    std_logic;
             DES_BUFFER_FREE : In    std_logic;
             DES_DATA_READY : In    std_logic;
             DES_ERR : In    std_logic;
             DES_PARITY : In    std_logic;
             DOUT_EMPTY : In    std_logic;
	     EQUAL : In    std_logic;
	     RESET : In    std_logic;
             RSA_NEXTEXP : In    std_logic;
             RSA_READY : In    std_logic;
             BUSY : Out   std_logic;
             DES_BUFFER_FREE_SET : Out   std_logic;
             DES_DATA_IS_KEY : Out   std_logic;
             DES_DATA_READY_SET : Out   std_logic;
             DES_IN_EN : Out   std_logic;
             DES_MODE : Out   std_logic_vector (4 downto 0);
             DEST_REG : Out   std_logic_vector (2 downto 0);
             ENABLE_TEST : Out   std_logic;
             EQ_REG : Out   std_logic;
             INT : Out   std_logic;
             RAM_SEL : Out   std_logic;
             RSA_GO : Out   std_logic;
             RSA_SEL : Out   std_logic_vector (1 downto 0);
             RSA_VAL_ACC : Out   std_logic;
             SOURCE_REG : Out   std_logic_vector (2 downto 0);
             STATE_EN : Out   std_logic;
             STATUS : Out   std_logic_vector (7 downto 0);
	     RAM_MODE : Out STD_LOGIC_VECTOR(5 downto 0);
	     RAM_ADR_IS_AT_END_OFF_ALL : In   std_logic;
	     RAM_ADR_IS_AT_END_OFF_TEMPEXP : In   std_logic;
	     RAM_ADR_IS_AT_END_OFF_MODUL : In   std_logic;
	     RAM_ADR_IS_AT_END_OFF_PUBLICKEY : In   std_logic;
	     RAM_ADR_IS_AT_END_OFF_PRIVATKEY : In   std_logic;
	     RAM_ADR_IS_AT_END_OFF_ZERTPUB : In   std_logic;
	     RAM_ADR_IS_AT_END_OFF_ZERTMODUL : In   std_logic;
	     INVERT : out std_logic );
end FSM_CORE;

architecture BEHAVIORAL of FSM_CORE is
    
    constant RSA_SEL_MODULO	: STD_LOGIC_VECTOR(1 downto 0) := "00";
    constant RSA_SEL_DATA	: STD_LOGIC_VECTOR(1 downto 0) := "01";
    constant RSA_SEL_KEY	: STD_LOGIC_VECTOR(1 downto 0) := "10";
    constant RSA_SEL_READ	: STD_LOGIC_VECTOR(1 downto 0) := "11";
    
    constant SEL_NOP		: STD_LOGIC_VECTOR(2 downto 0) := "000";
    constant SEL_LFSR_CONST	: STD_LOGIC_VECTOR(2 downto 0) := "000";  -- readonly
    constant SEL_IO		: STD_LOGIC_VECTOR(2 downto 0) := "001";
    constant SEL_RAM		: STD_LOGIC_VECTOR(2 downto 0) := "010";
    constant SEL_DES_LOW	: STD_LOGIC_VECTOR(2 downto 0) := "011";
    constant SEL_DES_HIGH	: STD_LOGIC_VECTOR(2 downto 0) := "100";
    constant SEL_RSA		: STD_LOGIC_VECTOR(2 downto 0) := "101";
    constant SEL_LFSR_LOW	: STD_LOGIC_VECTOR(2 downto 0) := "110";
    constant SEL_LFSR_HIGH	: STD_LOGIC_VECTOR(2 downto 0) := "111";
    
    type STATES is
	(
	    -- R E S E T 12
	    S_RESET,
	    S_DELETERAM,S_DELETERAM_END,
	    S_LOADRAM_BEGIN,S_LOADRAM_WAIT,S_LOADRAM_COPY,S_LOADRAM_END,
	    S_LOADFSM_WAIT1,S_LOADFSM_COPY1,S_LOADFSM_WAIT2,S_LOADFSM_COPY2,
	    S_PROTECT_CHIP,
	    -- C A R D C H A N G E 12
	    S_CARDCHANGE,
	    S_LOADPIN,S_LOADPIN_RAMACCESS,
	    S_WAITPIN,S_CHECKPIN_DECIDE,S_CHECKPIN_JUMP,
	    S_WAITPIN2,S_CHECKPIN_DECIDE2,S_CHECKPIN_JUMP2,
	    S_WAITPIN3,S_CHECKPIN_DECIDE3,S_CHECKPIN_JUMP3,
	    
	    -- N E W C O M M A N D 19
	    S_NEWCOMMAND,
	    S_ENCRYPT_RSA,S_RSA_KEY_WAIT,S_RSA_KEY_COPY,S_RSA_KEY_END,
	    S_RSA_MODULO_BEGIN,S_RSA_MODULO_WAIT,S_RSA_MODULO_COPY,S_RSA_MODULO_WAIT2,S_RSA_MODULO_END,
	    S_RSA_DATA_BEGIN,S_RSA_DATA_WAIT,S_RSA_DATA_COPY,S_RSA_DATA_WAIT2,S_RSA_DATA_END,
	    S_RSA_GO,S_RSA_SEL_TEMPEXP,S_RSA_SEL_PRIVATKEY,S_RSA_SEL_ZERTPUP,
	    
	    -- 13
	    S_RSA_EXP_WAIT,S_RSA_EXP_COPY,S_RSA_EXP_COPY_RAMACCESS,S_RSA_EXP_NEXT,
	    S_RSA_EXP_WAIT2,S_RSA_EXP_END,S_RSA_WAIT,
	    S_RSA_READ_BEGIN,S_RSA_READ_WAIT,S_RSA_READ_WAIT2,S_RSA_READ_COPY,S_RSA_READ_NEXT,S_RSA_READ_END,

	    -- 6
	    S_DECRYPT_RSA,S_DECRYPT_RSA_WAIT,S_DECRYPT_RSA_WRITE,S_DECRYPT_RSA_WRITE_RAMACCESS,
	    S_DECRYPT_RSA_COPY,S_DECRYPT_RSA_END,

	    -- 21
	    S_RSA2DES1_WAIT1,S_RSA2DES1_WAIT1B,S_RSA2DES1_WORD1,
	    S_RSA2DES1_WAIT2,S_RSA2DES1_WORD2, S_RSA2DES1_WAIT3, S_RSA2DES1_WRITE_KEY,
	    S_RSA2DES2_WAIT1,S_RSA2DES2_WAIT1B,S_RSA2DES2_WORD1,
	    S_RSA2DES2_WAIT2,S_RSA2DES2_WORD2, S_RSA2DES2_WAIT3, S_RSA2DES2_WRITE_KEY,
	    S_RSA2DES3_WAIT1,S_RSA2DES3_WAIT1B,S_RSA2DES3_WORD1,
	    S_RSA2DES3_WAIT2,S_RSA2DES3_WORD2, S_RSA2DES3_WAIT3, S_RSA2DES3_WRITE_KEY,

	    -- D E S  18
	    S_ENCRYPT_DES,S_DES_KEY1_GET1,S_DES_KEY1_WAIT,S_DES_KEY1_GET2,S_DES_KEY1_WAIT2,S_DES_KEY1_WRITE,
	    S_DES_KEY2,   S_DES_KEY2_GET1,S_DES_KEY2_WAIT,S_DES_KEY2_GET2,S_DES_KEY2_WAIT2,S_DES_KEY2_WRITE,
	    S_DES_KEY3,   S_DES_KEY3_GET1,S_DES_KEY3_WAIT,S_DES_KEY3_GET2,S_DES_KEY3_WAIT2,S_DES_KEY3_WRITE,

	    -- 10
	    S_DECRYPT_DES,

	    S_DES_READ_WRITE,
	    S_DES_WRITE_REG1,S_DES_WRITE_WAIT,S_DES_WRITE_REG2,S_DES_WRITE,
	    S_DES_READ_REG1,S_DES_READ_WAIT,S_DES_READ_REG2,S_DES_READ,

	    -- 23
	    S_MAKE_SIGNAUTURE,S_MAKE_SIG_INIT,S_MAKE_SIG_INIT2,
	    S_MAKE_SIG_WAIT1,S_MAKE_SIG_WAIT1A,S_MAKE_SIG_WAIT1B,
	    S_MAKE_SIG_WRITE1A,S_MAKE_SIG_WRITE1,S_MAKE_SIG_WAIT2,S_MAKE_SIG_WRITE2,S_MAKE_SIG_WRITE,
	    S_MAKE_SIG_RSA_WAIT1,S_MAKE_SIG_RSA_IGNORE,S_MAKE_SIG_RSA_COPY1,S_MAKE_SIG_RSA_WRITE1,
	    S_MAKE_SIG_RSA_WAIT2,S_MAKE_SIG_RSA_COPY2,S_MAKE_SIG_RSA_WRITE2,
	    S_MAKE_SIG_RSA_WAIT3,
	    S_MAKE_SIG_RSA_LFSR_COPY,S_MAKE_SIG_RSA_LFSR_WRITE,S_MAKE_SIG_RSA_LFSR_WAIT,S_MAKE_SIG_RSA_COPY4,

	    -- 2
	    S_AUTHENTIFY,
	    S_AUTHENTIFY_WAIT,

	    -- 22
	    S_CHECK_SIGNATURE,
	    S_CHECKSIGN_RSAREAD,S_CHECKSIGN_RSAREAD_COPY1,
	    S_CHECKSIGN_RSAREAD_WAIT2,S_CHECKSIGN_RSAREAD_COPY2,
	    S_CHECKSIGN_HASH,
	    S_CHECKSIGN_HASH_WAIT1B,S_CHECKSIGN_HASH_WRITE1,
	    S_CHECKSIGN_HASH_WAIT2, S_CHECKSIGN_HASH_WRITE2,
	    S_CHECKSIGN_HASH_WRITE,S_CHECKSIGN_HASH_WAIT3,
	    S_CHECKSIGN_HASH_NOKEY,
	    S_CHECKSIGN_ISEQ_LOW_LOAD,S_CHECKSIGN_ISEQ_LOW_CHECK_RAMACCESS,
	    S_CHECKSIGN_ISEQ_LOW_CHECK, S_CHECKSIGN_ISEQ_LOW_JUMP,
	    S_CHECKSIGN_ISEQ_HIGH_LOAD,S_CHECKSIGN_ISEQ_HIGH_CHECK_RAMACCESS,
	    S_CHECKSIGN_ISEQ_HIGH_CHECK, S_CHECKSIGN_ISEQ_HIGH_JUMP,
	    S_CHECKSIGN_ISEQ_OK,

	    -- 52
	    S_CHECK_AUTHENTIFY,S_CHECKAUTH_INIT,
	    S_CHECKAUTH_PREHASH_WAIT,
	    S_CHECKAUTH_PREHASH_COPY_L,
	    S_CHECKAUTH_PREHASH_COPY_H,
	    S_CHECKAUTH_PREHASH_WAIT2,
	    S_CHECKAUTH_PREHASH_COPYBACK_L,
	    S_CHECKAUTH_PREHASH_COPYBACK_H,
	    S_CHECKAUTH_OL_WAIT,S_CHECKAUTH_OL_COPY,S_CHECKAUTH_OH_WAIT_RAMACCESS,
	    S_CHECKAUTH_OH_WAIT,S_CHECKAUTH_OH_COPY,S_CHECKAUTH_HASH_WAIT_RAMACCESS,
	    S_CHECKAUTH_HASH_WAIT,S_CHECKAUTH_HASH_COPY_L,
	    S_CHECKAUTH_HASH_COPY_H,S_CHECKAUTH_HASH_COPY_H_RAMACCESS,
	    S_CHECKAUTH_HASH_WAIT2,S_CHECKAUTH_HASH_WAIT2_RAMACCESS,
	    S_CHECKAUTH_HASH_COPYBACK_L,S_CHECKAUTH_HASH_COPYBACK_H,	    
	    S_CHECKAUTH_RRSA_WAIT1,S_CHECKAUTH_RRSA_WORD1,
	    S_CHECKAUTH_RRSA_CHECK,S_CHECKAUTH_RRSA_CHECK_RAMACCESS,S_CHECKAUTH_RRSA_WAIT2,
	    S_CHECKAUTH_RRSA_WAIT2B,S_CHECKAUTH_RRSA_WORD2,S_CHECKAUTH_RRSA_DECIDE,
	    S_CHECKAUTH_RRSA_DECIDE_RAMACCESS,S_CHECKAUTH_RRSA_JUMP,S_CHECKAUTH_OK,
	    S_CHECKAUTH_HASH2_COPY_L_RAMACCESS,S_CHECKAUTH_HASH2_COPY_L,
	    S_CHECKAUTH_HASH2_COPY_H_RAMACCESS,S_CHECKAUTH_HASH2_COPY_H,
	    S_CHECKAUTH_HASH2_WAIT,
	    S_CHECKAUTH_HASH2_COPY2_L_RAMACCESS,S_CHECKAUTH_HASH2_COPY2_L,
	    S_CHECKAUTH_HASH2_COPY2_H_RAMACCESS,S_CHECKAUTH_HASH2_COPY2_H,
	    S_CHECKAUTH_HASH2_WAIT2,
	    S_CHECKAUTH_HASH2_IGNORE,
	    S_CHECKAUTH_HASH2_COPYBACK,S_CHECKAUTH_HASH2_COPYBACK_L,S_CHECKAUTH_HASH2_COPYBACK_H,	    
	    S_CHECKAUTH_RSA_MODUL_COPY,S_CHECKAUTH_RSA_MODUL_COPY_RAMACCESS,
	    S_CHECKAUTH_RSA_MODUL_WRITE,S_CHECKAUTH_RSA_MODUL_WAIT,
	    S_CHECKAUTH_OK2,

	    -- 6
	    S_SET_PIN,S_SET_PIN_LOAD,

	    S_SET_ZERT,S_SET_ZERT_WAIT,S_SET_ZERT_COPY,S_SET_ZERT_END,

	    -- 24
	    S_READ_PUBLIC_KEYS, S_READ_PUBLIC_KEYS_WAIT,
	    S_READ_PUBLIC_KEYS_COPY,S_READ_PUBLIC_KEYS_COPY_RAMACCESS,
	    S_READ_PUBLIC_KEYS_NEXT, S_READ_PUBLIC_KEYS_END, S_READ_PUBLIC_KEYS_NEXT2,

	    S_READ_USER_DATA, S_READ_USER_DATA_WAIT,
	    S_READ_USER_DATA_COPY,S_READ_USER_DATA_COPY_RAMACCES,
	    S_READ_USER_DATA_NEXT, S_READ_USER_DATA_END,

	    S_NAME_OUT, S_NAME_OUT_COPY, S_NAME_OUT_NEXT,

	    S_RAMTEST_WAIT_EXPECTED,S_RAMTEST_COPY_EXPECTED,
	    S_RAMTEST_WAIT_DATA,S_RAMTEST_CHECK,
	    S_RAMTEST_WRITE,S_RAMTEST_FAIL,S_RAMTEST_NEXT,
	    
	    S_IDLE
	);

    attribute enum_encoding : string;
    attribute enum_encoding of STATES: type is
	"0000000000000000000000 "&  	-- S_RESET
        "0000000100000101101111 "&
	"0000001000000000001111 "&
	"0000001100000000001111 "&
	"0000010000000000001111 "&
	"0000010100000100011111 "&
	"0000011000000000001111 "&
	"0000011100000000001111 "&
	"0000100000001110011111 "&
	"0000100100001100001111 "&
	"0000101000001100011111 "&
	"0000101100000000000111 "&  	-- S_PROTECT_CHIP
	"0000110000000000000111 "&  	-- S_CARDCHANGE
	"0000110100000000101111 "&
	"0000111001000000101111 "&
	"0000111100000000001111 "&
	"0001000000000000011111 "&
	"0001000100000000001111 "&
	"0001001000000000001111 "&
	"0001001100000000011111 "&
	"0001010000000000001111 "&
	"0001010100000000001111 "&
	"0001011000000000011111 "&
	"0001011100000000001111 "&  	-- S_CHECKPIN_JUMP3
	"0001100000000000001111 "&  	-- S_NEWCOMMAND
	"0001100100000000001111 "&
	"0001101000000000001111 "&
	"0001101100000100011111 "&
	"0001110000000000001111 "&
	"0001110100000000001001 "&
	"0001111000000000001111 "&
	"0001111100001010011111 "&
	"0010000000010000001111 "&
	"0010000100000000001111 "&
	"0010001000000000001101 "&
	"0010001100000000001111 "&
	"0010010000001010011111 "&
	"0010010100010000001111 "&
	"0010011000000000001111 "&
	"0010011100100000001011 "&
	"0010100000000000001111 "&
	"0010100100000000001111 "&
	"0010101000000000001111 "&  	-- S_RSA_SEL_ZERTPUP 
	"0010101100000000001111 "&  	-- S_RSA_EXP_WAIT
	"0010110000001010101111 "&
	"0010110100001010101111 "&
	"0010111000000000001111 "&
	"0010111100010000001111 "&
	"0011000000000000001111 "&
	"0011000100000000001111 "&
	"0011001000000000001111 "&
	"0011001100000000001111 "&
	"0011010000000000001111 "&
	"0011010100000011011111 "&
	"0011011000000000001111 "&
	"0011011100010000001111 "&  	-- S_RSA_READ_END
	"1111101100001000011111 "&      -- S_DECRYPT_RSA ----------------------
	"0011100000000000001001 "&  	-- S_DECRYPT_RSA_WAIT
	"0011100100000000001111 "&
	"0011101000010000001111 "&
	"0011101100001010101111 "&
	"0011110000000000101111 "&  	-- S_DECRYPT_RSA_END
	"0011110100000000001111 "&	-- S_RSA2DES1_WAIT1
	"0011111000000000001111 "&
	"0011111100000000001111 "&
	"0100000000010111011111 "&
	"0100000100000000001111 "&
	"0100001000011001011111 "&
	"0100001100000000001111 "&
	"0100010000000000001111 "&
	"0100010100000000001111 "&
	"0100011000000000001111 "&
	"0100011100010111011111 "&
	"0100100000000000001111 "&
	"0100100100011001011111 "&
	"0100101000000000001111 "&
	"0100101100000000001111 "&
	"0100110000000000001111 "&
	"0100110100000000001111 "&
	"0100111000010111011111 "&
	"0100111100000000001111 "&
	"0101000000011001011111 "&	-- S_RSA2DES3_WAIT3
	"1111110000000000001111 "&	-- S_RSA2DES3_WRITE_KEY ---------------
	"0101000100000000001111 "&	-- S_ENCRYPT_DES
	"0101001000000000001111 "&
	"0101001100000000001111 "&
	"0101010000000110011111 "&
	"0101010100000000001111 "&
	"0101011000001000011111 "&
	"0101011100000000001111 "&
	"0101100000000000001111 "&
	"0101100100000000001111 "&
	"0101101000000110011111 "&
	"0101101100000000001111 "&
	"0101110000001000011111 "&
	"0101110100000000001111 "&
	"0101111000000000001111 "&
	"0101111100000000001111 "&
	"0110000000000110011111 "&  	-- S_DES_KEY3_GET
	"1111110100000000001111 "&  	-- S_DES_KEY3_WAIT2 -------------------
	"0110000100000000001111 "&	-- S_DES_KEY3_WRITE
	"0110001000001000011111 "&
	"0110001100000000001111 "&
	"0110010000000000001111 "&
	"0110010100000000001001 "&
	"0110011000000000001110 "&
	"0110011100000110011111 "&
	"0110100000000000001111 "&
	"0110100100001000011111 "&
	"0110101000000000001111 "&
	"0110101100000010111111 "&  	-- S_DES_READ
	"0110110000000000001111 "&  	-- S_MAKE_SIGNAUTURE
	"0110110100000011001111 "&  	-- S_MAKE_SIG_INIT
	"1111111000000000001111 "&  	-- S_MAKE_SIG_INIT2--------------------
	"0110111000000000001111 "&  	-- S_MAKE_SIG_WAIT1
	"0110111100000010001111 "&
	"0111000000000000001111 "&
	"0111000100000000001111 "&
	"0111001000000000001111 "&
	"0111001100000000001111 "&
	"0111010000000000001111 "&
	"0111010100000110011111 "&
	"0111011000000110011110 "&
	"0111011100000000001111 "&
	"0111100000001000011111 "&
	"0111100100000000001111 "&
	"0111101000000000001101 "&
	"0111101100000000001111 "&
	"0111110000001010111111 "&
	"0111110100010000001111 "&
	"0111111000000000001111 "&
	"0111111100001011001111 "&
	"1000000000010000001111 "&
	"1000000100000000001111 "&  	-- S_MAKE_SIG_RSA_COPY4
	"1000001000001011101111 "&  	-- S_AUTHENTIFY
	"1000001100010000001111 "&	-- S_AUTHENTIFY_WAIT
	"1000010000000000001111 "&  	-- S_CHECK_SIGNATURE
	"1000010100011010001111 "&
	"1000011000000000001111 "&
	"1000011100000000001111 "&
	"1000100000000000001111 "&
	"1000100100000011101111 "&
	"1000101000010101011111 "&
	"1000101100000000001111 "&
	"1000110000010101011111 "&
	"1000110100000000001111 "&
	"1000111000000000001111 "&
	"1000111100000110011111 "&
	"1001000000000000001111 "&
	"1001000100001000011111 "&
	"1001001000000000001111 "&
	"1001001100000000001111 "&
	"1001010000000000001110 "&
	"1001010100000000101110 "&
	"1001011001000000101111 "&
	"1001011100000000111111 "&
	"1001100000000000001111 "&
	"1001100101000000101111 "&  	-- S_CHECKSIGN_ISEQ_OK
	"1001101001000000101111 "&  	-- S_CHECK_AUTHENTIFY
	"1111111100000000001111 "&  	-- S_CHECKAUTH_INIT -------------------
	"1001101100000001001111 "&  	-- S_CHECKAUTH_PREHASH_WAIT
	"1001110000000000001111 "&
	"1001110100000000001111 "&
	"1001111000000000001111 "&
	"1001111100000000001111 "&
	"1010000000000000001111 "&
	"1010000100000111101111 "&
	"1010001000001001111111 "&
	"1010001100000000001111 "&
	"1010010000000100111111 "&
	"1010010100000101001111 "&
	"1010011000000000001111 "&
	"1010011100000000101111 "&
	"1010100000000010101111 "&
	"1010100100000000001111 "&
     	"1010101000000000101111 "&
	"1010101100000010101111 "&
	"1010110000000000001111 "&
	"1010110100000000101111 "&
	"1010111000000000101111 "&
	"1010111100000110101111 "&
	"1011000000000000001111 "&
	"1011000100001000101111 "&
	"1011001000000100111111 "&
	"1011001100000101001111 "&
	"1011010000000000001111 "&
	"1011010101000001011111 "&
	"1011011000000000101111 "&
	"1011011100000000101111 "&
	"1011100000010000001111 "&
	"1011100100000000001111 "&
	"1011101001010001011111 "&
	"1011101100000000101111 "&
	"1011110000000000101111 "&
	"1011110100000000001111 "&
	"1011111000000000001111 "&
	"1011111100000110101111 "&
	"1100000000000000101111 "&
	"1100000100001000101111 "&
	"1100001000000000101111 "&
	"1100001100000000001111 "&
	"1100010000000110101111 "&
	"1100010100000000101111 "&
	"1100011000001000101110 "&
	"1100011100000000101111 "&
	"1100100000000000001111 "&
	"1100100100000000001111 "&
	"1100101000000000001111 "&
	"1100101100000100111111 "&
	"1100110000000101001001 "&  	-- S_CHECKAUTH_OK2
	"1100110100000000101111 "&  	-- S_SET_PIN
	"1100111000001010101111 "&
	"1100111100010000001111 "&
	"1101000000000000001111 "&
	"1101000100000000000111 "&
	"1101001000000000001111 "&  	-- S_SET_ZERT_END
	"1101001100000100011111 "&  	-- S_READ_PUBLIC_KEYS
	"1101010000000000001111 "&
	"1101010100000000001111 "&
	"1101011000000100011111 "&
	"1101011100000000001111 "&
	"1101100000000000001111 "&
	"1101100100000000001111 "&
	"1101101000000000101111 "&
	"1101101100000010101111 "&
	"1101110000000000001111 "&
	"1101110100000000001111 "&
	"1101111000000000001111 "&
	"1101111100000000001111 "&
	"1110000000000000001111 "&
	"1110000100000000101111 "&
	"1110001000000010101111 "&
	"1110001100000000001111 "&
	"1110010000000000001111 "&
	"1110010110000000001111 "&
	"1110011010000010101111 "&
	"1110011110000000001111 "&
	"1110100000000000001111 "&
	"1110100101000000011111 "&
	"1110101000000000101111 ";  	-- S_IDLE

    signal NEWSTATE : STATES;
    signal STATE : STATES;
    attribute state_vector : string;
    attribute state_vector of BEHAVIORAL : architecture is "STATE";

    subtype SECURITY_LEVEL is STD_LOGIC_VECTOR(1 downto 0);
    constant NO_KEY		: SECURITY_LEVEL := "00";
    constant SECRET_KEY		: SECURITY_LEVEL := "01";
    constant AUTHENTIFIED	: SECURITY_LEVEL := "10";
    constant SPECIAL_MODE	: SECURITY_LEVEL := "11";
    signal SECURITY : SECURITY_LEVEL;
    signal OLD_SECURITY : SECURITY_LEVEL;

    signal RESULT_I : STD_LOGIC;
    signal OLD_RESULT_I : STD_LOGIC;

    signal RSA_SEL_I : STD_LOGIC_VECTOR(1 downto 0);
    signal OLD_RSA_SEL_I : STD_LOGIC_VECTOR(1 downto 0);

    signal DES_DATA_IS_KEY_I : STD_LOGIC;
    signal OLD_DES_DATA_IS_KEY_I : STD_LOGIC;

begin
    
    -- purpose: speicherung des zustands, reset
    process(CLK,RESET)
    begin
	if RESET='1' then
	    STATE <= S_RESET;
	    OLD_SECURITY <= SECRET_KEY;
	    OLD_RESULT_I <= '0';
	    OLD_RSA_SEL_I <= RSA_SEL_MODULO;
	    OLD_DES_DATA_IS_KEY_I <= '1';
	elsif CLK'event AND CLK='1' then
	    if CARDCHANGE='0' and STATE >= S_NEWCOMMAND then -- for more security
		STATE <= S_CARDCHANGE;
	    elsif CTRL_CHANGE='1'
	      and ( (STATE >= S_NEWCOMMAND)
	       or   (SECURITY = NO_KEY) ) then -- for more security
		STATE <= S_NEWCOMMAND;
	    else
		STATE <= NEWSTATE;
	    end if;
	    OLD_SECURITY <= SECURITY;
	    OLD_RESULT_I <= RESULT_I;
	    OLD_RSA_SEL_I <= RSA_SEL_I;
	    OLD_DES_DATA_IS_KEY_I <= DES_DATA_IS_KEY_I;
	end if;
    end process;

    
    process(STATE, CTRL, DATA_VALID, DES_ERR, DES_PARITY, DOUT_EMPTY,DES_BUFFER_FREE,
	   DES_DATA_READY, EQUAL, RSA_NEXTEXP, RSA_READY, SECURITY, RESULT_I,
	   RAM_ADR_IS_AT_END_OFF_ALL, RAM_ADR_IS_AT_END_OFF_TEMPEXP,
	   RAM_ADR_IS_AT_END_OFF_MODUL, RAM_ADR_IS_AT_END_OFF_PUBLICKEY,
	   RAM_ADR_IS_AT_END_OFF_PRIVATKEY, RAM_ADR_IS_AT_END_OFF_ZERTPUB,
	   RAM_ADR_IS_AT_END_OFF_ZERTMODUL,
	   OLD_DES_DATA_IS_KEY_I, OLD_RSA_SEL_I, OLD_RESULT_I, OLD_SECURITY )
    begin
        SECURITY <= OLD_SECURITY;
        RESULT_I <= OLD_RESULT_I;
        RSA_SEL_I <= OLD_RSA_SEL_I;
        DES_DATA_IS_KEY_I  <= OLD_DES_DATA_IS_KEY_I;
	NEWSTATE <= S_RESET;
	DES_DATA_READY_SET <= '0';
	DES_BUFFER_FREE_SET <= '0';
	DEST_REG <= "000";
	EQ_REG <= '0';
	BUSY <= '0';
        RAM_MODE <= RAM_MODE_NOP;
	RSA_GO <= '0';
        RSA_VAL_ACC <='0';
	SOURCE_REG <= "000";
	STATE_EN <= '1'; -- fest ?
        RAM_SEL <= '0';

	case STATE is
	    -- reset --
	    when S_RESET =>
		RSA_SEL_I	<= RSA_SEL_MODULO;
	        SECURITY <= SECRET_KEY;
		RAM_MODE <= RAM_MODE_SET_PUBLICKEY;
		DES_BUFFER_FREE_SET <= '1';
		DES_DATA_IS_KEY_I <= '0';
		NEWSTATE <= S_DELETERAM;

	    when S_DELETERAM =>
		SOURCE_REG <= SEL_LFSR_LOW;
		DEST_REG <= SEL_RAM;
		RAM_MODE <= RAM_MODE_INC;
		NEWSTATE <= S_DELETERAM_END;
	    when S_DELETERAM_END =>
		if RAM_ADR_IS_AT_END_OFF_ALL /= '1' then
		    NEWSTATE <= S_DELETERAM;
		else
		    NEWSTATE <= S_LOADRAM_BEGIN;
		end if;
		
	    when S_LOADRAM_BEGIN =>
		SECURITY <= NO_KEY;
		RAM_MODE <= RAM_MODE_SET_PUBLICKEY;
		NEWSTATE <= S_LOADRAM_WAIT;
	    when S_LOADRAM_WAIT =>
		if DATA_VALID='1' then
		    NEWSTATE <= S_LOADRAM_COPY;
		else
		    NEWSTATE <= S_LOADRAM_WAIT;
		end if;
	    when S_LOADRAM_COPY =>
		SOURCE_REG <= SEL_IO;
		DEST_REG <= SEL_RAM;
		RAM_MODE <= RAM_MODE_INC;
		NEWSTATE <= S_LOADRAM_END;
	    when S_LOADRAM_END =>
		if RAM_ADR_IS_AT_END_OFF_ALL /= '1' then
		    NEWSTATE <= S_LOADRAM_WAIT;
		else
		    NEWSTATE <= S_LOADFSM_WAIT1;
		end if;
		
	    when S_LOADFSM_WAIT1 =>
		if DATA_VALID='1' then
		    NEWSTATE <= S_LOADFSM_COPY1;
		else
		    NEWSTATE <= S_LOADFSM_WAIT1;
		end if;
	    when S_LOADFSM_COPY1 =>
		SOURCE_REG <= SEL_IO;
		DEST_REG <= SEL_LFSR_HIGH;
		NEWSTATE <= S_LOADFSM_WAIT2;
	    when S_LOADFSM_WAIT2 =>
		DEST_REG <= SEL_LFSR_LOW;
		if DATA_VALID='1' then
		    NEWSTATE <= S_LOADFSM_COPY2;
		else
		    NEWSTATE <= S_LOADFSM_WAIT2;
		end if;
	    when S_LOADFSM_COPY2 =>
		BUSY <= '1';
		SOURCE_REG <= SEL_IO;
		DEST_REG <= SEL_LFSR_LOW;
		NEWSTATE <= S_PROTECT_CHIP;
		
	    when S_PROTECT_CHIP =>
		BUSY <= '1';
		SECURITY <= AUTHENTIFIED;
		NEWSTATE <= S_IDLE;

	    -- card-change (enter pin 3 try's else delete keys)--
	    when S_CARDCHANGE =>
		BUSY <= '1';
		SECURITY <= SECRET_KEY;
		RAM_MODE <= RAM_MODE_SET_PIN;
		NEWSTATE <= S_LOADPIN;
	    when S_LOADPIN =>
		SOURCE_REG <= SEL_RAM;  --1
		NEWSTATE <= S_LOADPIN_RAMACCESS;
	    when S_LOADPIN_RAMACCESS =>
		SOURCE_REG <= SEL_RAM;  --2
		EQ_REG <= '1';
      		if DATA_VALID='1' then
		    NEWSTATE <= S_CHECKPIN_DECIDE;
		else
		    NEWSTATE <= S_WAITPIN;
		end if;

	    when S_WAITPIN =>
      		if DATA_VALID='1' then
		    NEWSTATE <= S_CHECKPIN_DECIDE;
		else
		    NEWSTATE <= S_WAITPIN;
		end if;		
	    when S_CHECKPIN_DECIDE =>
		SOURCE_REG <= SEL_IO;
		NEWSTATE <= S_CHECKPIN_JUMP;
	    when S_CHECKPIN_JUMP =>
		if EQUAL = '1' then
		    NEWSTATE <= S_IDLE;
		else 
		    NEWSTATE <= S_WAITPIN2;
		end if;

	    when S_WAITPIN2 =>  	-- two tries left
      		if DATA_VALID='1' then
		    NEWSTATE <= S_CHECKPIN_DECIDE2;
		else
		    NEWSTATE <= S_WAITPIN2;
		end if;
	    when S_CHECKPIN_DECIDE2 =>	
		SOURCE_REG <= SEL_IO;
		NEWSTATE <= S_CHECKPIN_JUMP2;
	    when S_CHECKPIN_JUMP2 =>
		if EQUAL = '1' then
		    NEWSTATE <= S_IDLE;
		else 
		    NEWSTATE <= S_WAITPIN3;
		end if;
		
	    when S_WAITPIN3 =>  	-- last change
      		if DATA_VALID='1' then
		    NEWSTATE <= S_CHECKPIN_DECIDE3;
		else
		    NEWSTATE <= S_WAITPIN3;
		end if;
	    when S_CHECKPIN_DECIDE3 =>
		SOURCE_REG <= SEL_IO;
		NEWSTATE <= S_CHECKPIN_JUMP3;
	    when S_CHECKPIN_JUMP3 =>
		if EQUAL = '1' then
		    NEWSTATE <= S_IDLE;
		else 
		    NEWSTATE <= S_RESET;
		end if;
		
	    -- new-command --
	    when S_NEWCOMMAND =>
		RAM_MODE <= RAM_MODE_SET_PUBLICKEY;
		DES_BUFFER_FREE_SET <= '1';
		
		NEWSTATE <= S_IDLE;
		
		case CTRL(4 downto 0) is
		    when "00001" =>
			NEWSTATE <= S_ENCRYPT_RSA;
		    when "01001" =>
			NEWSTATE <= S_DECRYPT_RSA;
		    when "10000"|"10001"|"10010"|"10011"|"10100"|"10101"|"10110"|"10111" =>
			NEWSTATE <= S_ENCRYPT_DES;
		    when "11000"|"11001"|"11010"|"11011"|"11100"|"11101"|"11110"|"11111" =>
			NEWSTATE <= S_DECRYPT_DES;
		    when "01011" =>
			NEWSTATE <= S_MAKE_SIGNAUTURE;
		    when "00011" =>
			NEWSTATE <= S_CHECK_SIGNATURE;
		    when "00010" =>
			NEWSTATE <= S_AUTHENTIFY;
		    when "00000" =>
			NEWSTATE <= S_CHECK_AUTHENTIFY;
		    when "01100" =>
			NEWSTATE <= S_SET_PIN;
		    when "01101" =>
			NEWSTATE <= S_SET_ZERT;
		    when "00110" =>
			NEWSTATE <= S_READ_PUBLIC_KEYS;
		    when "01111" =>
			NEWSTATE <= S_READ_USER_DATA;
		    when "01000" =>
			NEWSTATE <= S_NAME_OUT;
		    when others =>
			NEWSTATE <= S_IDLE;
		end case;
		
		if (CTRL(4 downto 0) = "01010") and (SECURITY = NO_KEY) then
		    NEWSTATE <= S_RAMTEST_WAIT_EXPECTED;
		elsif (CTRL(4 downto 3) = "11") and (SECURITY = NO_KEY) then
		    NEWSTATE <= S_ENCRYPT_DES;
		elsif CTRL(3) = '1' and SECURITY /= AUTHENTIFIED then
		    NEWSTATE <= S_IDLE;
		end if;

	    when S_ENCRYPT_RSA =>  	-- copy key to ram
		RAM_MODE <= RAM_MODE_SET_TEMPEXP;
		NEWSTATE <= S_RSA_KEY_WAIT;
	    when S_RSA_KEY_WAIT =>
		if DATA_VALID = '1' then
		    NEWSTATE <= S_RSA_KEY_COPY;
		else
		    NEWSTATE <= S_RSA_KEY_WAIT;
		end if;
	    when S_RSA_KEY_COPY =>
		SOURCE_REG <= SEL_IO;
		DEST_REG <= SEL_RAM;
		RAM_MODE <= RAM_MODE_INC;
		NEWSTATE <= S_RSA_KEY_END;
	    when S_RSA_KEY_END =>
		if RAM_ADR_IS_AT_END_OFF_TEMPEXP /= '1' then
		    NEWSTATE <= S_RSA_KEY_WAIT;
		else
		    NEWSTATE <= S_RSA_MODULO_BEGIN;
		end if;
		
	    when S_RSA_MODULO_BEGIN =>  -- move modulo from io to rsa
		RSA_SEL_I <= RSA_SEL_MODULO;
		RAM_MODE <= RAM_MODE_SET_MODUL;  -- counter
		NEWSTATE <= S_RSA_MODULO_WAIT;
	    when S_RSA_MODULO_WAIT =>
		if DATA_VALID = '1' then
		    NEWSTATE <= S_RSA_MODULO_COPY;
		else
		    NEWSTATE <= S_RSA_MODULO_WAIT;
		end if;
	    when S_RSA_MODULO_COPY =>
		SOURCE_REG <= SEL_IO;
		DEST_REG <= SEL_RSA;
		RAM_MODE <= RAM_MODE_INC;
		NEWSTATE <= S_RSA_MODULO_WAIT2;
	    when S_RSA_MODULO_WAIT2 =>
		RSA_VAL_ACC <= '1';
		if RSA_READY = '0' then
		    NEWSTATE <= S_RSA_MODULO_END;
		elsif RAM_ADR_IS_AT_END_OFF_MODUL /= '1' then
		    NEWSTATE <= S_RSA_MODULO_WAIT;
		else
		    NEWSTATE <= S_RSA_DATA_BEGIN;
		end if;
	    when S_RSA_MODULO_END =>
		if RSA_READY = '0' then
		    NEWSTATE <= S_RSA_MODULO_END;
		elsif RAM_ADR_IS_AT_END_OFF_MODUL /= '1' then
		    NEWSTATE <= S_RSA_MODULO_WAIT;
		else
		    NEWSTATE <= S_RSA_DATA_BEGIN;
		end if;

	    when S_RSA_DATA_BEGIN =>  	-- move data from io to rsa
		RSA_SEL_I <= RSA_SEL_DATA;
		RAM_MODE <= RAM_MODE_SET_PUBLICKEY;  -- counter
		NEWSTATE <= S_RSA_DATA_WAIT;
	    when S_RSA_DATA_WAIT =>
		if DATA_VALID = '1' then
		    NEWSTATE <= S_RSA_DATA_COPY;
		else
		    NEWSTATE <= S_RSA_DATA_WAIT;
		end if;
	    when S_RSA_DATA_COPY =>
		SOURCE_REG <= SEL_IO;
		DEST_REG <= SEL_RSA;
		RAM_MODE <= RAM_MODE_INC;
		NEWSTATE <= S_RSA_DATA_WAIT2;
	    when S_RSA_DATA_WAIT2 =>
		RSA_VAL_ACC <= '1';
		if RSA_READY = '0' then
		    NEWSTATE <= S_RSA_DATA_END;
		elsif RAM_ADR_IS_AT_END_OFF_PUBLICKEY /= '1' then
		    NEWSTATE <= S_RSA_DATA_WAIT;
		else
		    NEWSTATE <= S_RSA_GO;
	        end if;
	    when S_RSA_DATA_END =>
		if RSA_READY = '0' then
		    NEWSTATE <= S_RSA_DATA_END;
		elsif RAM_ADR_IS_AT_END_OFF_PUBLICKEY /= '1' then
		    NEWSTATE <= S_RSA_DATA_WAIT;
		else
		    NEWSTATE <= S_RSA_GO;
	        end if;

	    when S_RSA_GO =>
		RSA_GO <= '1';
		RSA_SEL_I <= RSA_SEL_KEY;
		if  CTRL(3) = '1'  -- secure Operation
		    and SECURITY = AUTHENTIFIED then
		    NEWSTATE <= S_RSA_SEL_PRIVATKEY;
		else
		    if CTRL(4 downto 0)="00000" and RESULT_I='1' then
			NEWSTATE <= S_RSA_SEL_ZERTPUP;
		    else
			NEWSTATE <= S_RSA_SEL_TEMPEXP;
		    end if;
		end if;
     	    when S_RSA_SEL_TEMPEXP =>
		RAM_MODE <= RAM_MODE_SET_TEMPEXP;
		NEWSTATE <= S_RSA_EXP_COPY;
     	    when S_RSA_SEL_ZERTPUP =>
		RAM_MODE <= RAM_MODE_SET_ZERTPUB;
		NEWSTATE <= S_RSA_EXP_COPY;
	    when S_RSA_SEL_PRIVATKEY =>
		RAM_MODE <= RAM_MODE_SET_PRIVATKEY;
		NEWSTATE <= S_RSA_EXP_COPY;
	    when S_RSA_EXP_COPY =>
		SOURCE_REG <= SEL_RAM;  --1
		DEST_REG <= SEL_RSA;
		NEWSTATE <= S_RSA_EXP_COPY_RAMACCESS;
	    when S_RSA_EXP_COPY_RAMACCESS =>
		SOURCE_REG <= SEL_RAM;  --2
		DEST_REG <= SEL_RSA;
		NEWSTATE <= S_RSA_EXP_WAIT;
	    when S_RSA_EXP_WAIT =>
		if RSA_NEXTEXP = '1' then
		    NEWSTATE <= S_RSA_EXP_WAIT2;
		else
		    NEWSTATE <= S_RSA_EXP_WAIT;
		end if;
	    when S_RSA_EXP_WAIT2 =>
		RSA_VAL_ACC <= '1';
		if RSA_NEXTEXP = '0' then
		    NEWSTATE <= S_RSA_EXP_NEXT;
		else
		    NEWSTATE <= S_RSA_EXP_WAIT2;
		end if;
	    when S_RSA_EXP_NEXT =>
		RAM_MODE <= RAM_MODE_INC;
		NEWSTATE <= S_RSA_EXP_END;
	    when S_RSA_EXP_END =>
		if	RAM_ADR_IS_AT_END_OFF_PRIVATKEY /= '1'
		    and RAM_ADR_IS_AT_END_OFF_TEMPEXP /= '1'
		    and RAM_ADR_IS_AT_END_OFF_ZERTPUB /= '1'
		then
		    NEWSTATE <= S_RSA_EXP_COPY;
		else
		    NEWSTATE <= S_RSA_WAIT;
	        end if;

	    when S_RSA_WAIT =>
		if CTRL(4 downto 3)="11" then -- DES
		    NEWSTATE <= S_RSA2DES1_WAIT1;
		elsif CTRL(4 downto 0) = "00000" then  -- check authendify
		    NEWSTATE <= S_CHECKAUTH_RRSA_WAIT1;
		elsif CTRL(4 downto 0)="00011" then  -- check sign
		    NEWSTATE <= S_CHECKSIGN_RSAREAD;
		else		    		    
		    NEWSTATE <= S_RSA_READ_BEGIN;
		end if;

	    when S_RSA_READ_BEGIN =>
		RSA_SEL_I <= RSA_SEL_READ;
		RAM_MODE <= RAM_MODE_SET_PUBLICKEY;  -- counter
		NEWSTATE <= S_RSA_READ_WAIT;
	    when S_RSA_READ_WAIT =>
		if  RSA_READY='1' then
		    if DOUT_EMPTY = '1' then
			NEWSTATE <= S_RSA_READ_COPY;
		    else
			NEWSTATE <= S_RSA_READ_WAIT2;
		    end if;
		else
		    NEWSTATE <= S_RSA_READ_WAIT;
		end if;
	    when S_RSA_READ_WAIT2 =>
		if DOUT_EMPTY = '1' then
		    NEWSTATE <= S_RSA_READ_COPY;
		else
		    NEWSTATE <= S_RSA_READ_WAIT2;
		end if;
	    when S_RSA_READ_COPY =>
		SOURCE_REG <= SEL_RSA;
		DEST_REG <= SEL_IO;
		NEWSTATE <= S_RSA_READ_NEXT;
	    when S_RSA_READ_NEXT =>
		RAM_MODE <= RAM_MODE_INC;
		NEWSTATE <= S_RSA_READ_END;
	    when S_RSA_READ_END =>
		RSA_VAL_ACC <= '1';
		if RAM_ADR_IS_AT_END_OFF_PUBLICKEY /= '1' then
		    NEWSTATE <= S_RSA_READ_WAIT;
		else
		    NEWSTATE <= S_RSA_DATA_BEGIN;
	        end if;
		    
	    when S_DECRYPT_RSA | S_DECRYPT_DES =>  	-- copy modul from ram to rsa
		RSA_SEL_I <= RSA_SEL_MODULO;
		RAM_MODE <= RAM_MODE_SET_MODUL;  -- counter
		NEWSTATE <= S_DECRYPT_RSA_COPY;
	    when S_DECRYPT_RSA_COPY =>
		SOURCE_REG <= SEL_RAM;  --1
		NEWSTATE <= S_DECRYPT_RSA_WRITE_RAMACCESS;
	    when S_DECRYPT_RSA_WRITE_RAMACCESS =>
		RAM_MODE <= RAM_MODE_INC;
		SOURCE_REG <= SEL_RAM;  --2
		DEST_REG <= SEL_RSA;
		NEWSTATE <= S_DECRYPT_RSA_WRITE;
	    when S_DECRYPT_RSA_WRITE =>
		RSA_VAL_ACC <= '1';		
		NEWSTATE <= S_DECRYPT_RSA_WAIT;
	    when S_DECRYPT_RSA_WAIT =>
		if RSA_READY = '0' then
		    NEWSTATE <= S_DECRYPT_RSA_WAIT;
		else
		    NEWSTATE <= S_DECRYPT_RSA_END;
		end if;
	    when S_DECRYPT_RSA_END =>
		if RAM_ADR_IS_AT_END_OFF_MODUL /= '1' then
		    NEWSTATE <= S_DECRYPT_RSA_COPY;
		else
		    if CTRL(4 downto 0) = "01001" then
			NEWSTATE <= S_RSA_DATA_BEGIN;  -- decrypt_rsa
		    else
			NEWSTATE <= S_RSA_GO;
		    end if;
		end if;

	    when S_RSA2DES1_WAIT1 =>  	-- copy DES-Key from RSA to DES
		RSA_SEL_I <= RSA_SEL_READ;
		if RSA_READY = '1' then
		    if DES_DATA_READY = '0' then
			NEWSTATE <= S_RSA2DES1_WORD1;
		    else
			NEWSTATE <= S_RSA2DES1_WAIT1B;
		    end if;
		else
		    NEWSTATE <= S_RSA2DES1_WAIT1;
		end if;
	    when S_RSA2DES1_WAIT1B =>
		if DES_DATA_READY = '0' then                                                                   
		    NEWSTATE <= S_RSA2DES1_WORD1;
		else
		    NEWSTATE <= S_RSA2DES1_WAIT1B;
		end if;
	    when S_RSA2DES1_WORD1 =>
	        RSA_VAL_ACC <= '1';
		SOURCE_REG <= SEL_RSA;
		DEST_REG <= SEL_DES_LOW;
		NEWSTATE <= S_RSA2DES1_WAIT2;
	    when S_RSA2DES1_WAIT2 =>
		if RSA_READY = '0' then
		    NEWSTATE <= S_RSA2DES1_WAIT2;
		else
		    NEWSTATE <= S_RSA2DES1_WORD2;
		end if;
	    when S_RSA2DES1_WORD2 =>
	        RSA_VAL_ACC <= '1';
		SOURCE_REG <= SEL_RSA;
		DEST_REG <= SEL_DES_HIGH;
		NEWSTATE <= S_RSA2DES1_WRITE_KEY;
	    when S_RSA2DES1_WRITE_KEY =>
		DES_DATA_IS_KEY_I <= '1';
		DES_DATA_READY_SET <= '1';
		NEWSTATE <= S_RSA2DES1_WAIT3;
	    when S_RSA2DES1_WAIT3 => 
		if DES_DATA_READY = '1' then
		    NEWSTATE <= S_RSA2DES1_WAIT3;
		else
		    if CTRL(1 downto 0) /= "00" then
			NEWSTATE <= S_RSA2DES2_WAIT1;
		    else
			NEWSTATE <= S_DES_READ_WRITE;
		    end if;
		end if;
	    when S_RSA2DES2_WAIT1 =>
		if RSA_READY = '1' then
		    if DES_DATA_READY = '0' then
			NEWSTATE <= S_RSA2DES2_WORD1;
		    else
			NEWSTATE <= S_RSA2DES2_WAIT1B;
		    end if;
		else
		    NEWSTATE <= S_RSA2DES2_WAIT1;
		end if;
	    when S_RSA2DES2_WAIT1B =>
		if DES_DATA_READY = '0' then                                                                   
		    NEWSTATE <= S_RSA2DES2_WORD1;
		else
		    NEWSTATE <= S_RSA2DES2_WAIT1B;
		end if;
	    when S_RSA2DES2_WORD1 =>
	        RSA_VAL_ACC <= '1';
		SOURCE_REG <= SEL_RSA;
		DEST_REG <= SEL_DES_LOW;
		NEWSTATE <= S_RSA2DES2_WAIT2;
	    when S_RSA2DES2_WAIT2 =>
		if RSA_READY = '0' then
		    NEWSTATE <= S_RSA2DES2_WAIT2;
		else
		    NEWSTATE <= S_RSA2DES2_WORD2;
		end if;
	    when S_RSA2DES2_WORD2 =>
	        RSA_VAL_ACC <= '1';
		SOURCE_REG <= SEL_RSA;
		DEST_REG <= SEL_DES_HIGH;
		NEWSTATE <= S_RSA2DES2_WRITE_KEY;
	    when S_RSA2DES2_WRITE_KEY =>
		DES_DATA_IS_KEY_I <= '1';
		DES_DATA_READY_SET <= '1';
		NEWSTATE <= S_RSA2DES2_WAIT3;
	    when S_RSA2DES2_WAIT3 => 
		if DES_DATA_READY = '1' then
		    NEWSTATE <= S_RSA2DES2_WAIT3;
		else
		    if CTRL(1 downto 0) /= "01" then
			NEWSTATE <= S_RSA2DES3_WAIT1;
		    else
			NEWSTATE <= S_DES_READ_WRITE;
		    end if;
		end if;
	    when S_RSA2DES3_WAIT1 =>
		if RSA_READY = '1' then
		    if DES_DATA_READY = '0' then
			NEWSTATE <= S_RSA2DES3_WORD1;
		    else
			NEWSTATE <= S_RSA2DES3_WAIT1B;
		    end if;
		else
		    NEWSTATE <= S_RSA2DES3_WAIT1;
		end if;
	    when S_RSA2DES3_WAIT1B =>
		if DES_DATA_READY = '0' then                                                                   
		    NEWSTATE <= S_RSA2DES3_WORD1;
		else
		    NEWSTATE <= S_RSA2DES3_WAIT1B;
		end if;
	    when S_RSA2DES3_WORD1 =>
	        RSA_VAL_ACC <= '1';
		SOURCE_REG <= SEL_RSA;
		DEST_REG <= SEL_DES_LOW;
		NEWSTATE <= S_RSA2DES3_WAIT2;
	    when S_RSA2DES3_WAIT2 =>
		if RSA_READY = '0' then
		    NEWSTATE <= S_RSA2DES3_WAIT2;
		else
		    NEWSTATE <= S_RSA2DES3_WORD2;
		end if;
	    when S_RSA2DES3_WORD2 =>
	        RSA_VAL_ACC <= '1';
		SOURCE_REG <= SEL_RSA;
		DEST_REG <= SEL_DES_HIGH;
		NEWSTATE <= S_RSA2DES3_WRITE_KEY;
	    when S_RSA2DES3_WRITE_KEY =>
		DES_DATA_IS_KEY_I <= '1';
		DES_DATA_READY_SET <= '1';
		NEWSTATE <= S_RSA2DES3_WAIT3;
	    when S_RSA2DES3_WAIT3 => 
		if DES_DATA_READY = '1' then
		    NEWSTATE <= S_RSA2DES3_WAIT3;
		else
		    NEWSTATE <= S_DES_READ_WRITE;
		end if;

	    when S_ENCRYPT_DES =>
		if DES_DATA_READY = '1' or DATA_VALID = '0' then
		    NEWSTATE <= S_ENCRYPT_DES;
		else
		    NEWSTATE <= S_DES_KEY1_GET1;
		end if;
	    when S_DES_KEY1_GET1 =>
		SOURCE_REG <= SEL_IO;
		DEST_REG <= SEL_DES_LOW;
		NEWSTATE <= S_DES_KEY1_WAIT;
	    when S_DES_KEY1_WAIT =>
		if DATA_VALID = '0' then
		    NEWSTATE <= S_DES_KEY1_WAIT;
		else
		    NEWSTATE <= S_DES_KEY1_GET2;
		end if;
	    when S_DES_KEY1_GET2 =>
		SOURCE_REG <= SEL_IO;
		DEST_REG <= SEL_DES_HIGH;
		NEWSTATE <= S_DES_KEY1_WRITE;				
	    when S_DES_KEY1_WRITE =>
		DES_DATA_IS_KEY_I <= '1';
		DES_DATA_READY_SET <= '1';
		NEWSTATE <= S_DES_KEY1_WAIT2;
	    when S_DES_KEY1_WAIT2 => 
		if DES_DATA_READY = '1' then
		    NEWSTATE <= S_DES_KEY1_WAIT2;
		else
		    if CTRL(1 downto 0) /= "00" then
			NEWSTATE <= S_DES_KEY2;
		    else
			NEWSTATE <= S_DES_READ_WRITE;
		    end if;
		end if;
	    when S_DES_KEY2 =>
		if DES_DATA_READY = '1' or DATA_VALID = '0' then
		    NEWSTATE <= S_DES_KEY2;
		else
		    NEWSTATE <= S_DES_KEY2_GET1;
		end if;
	    when S_DES_KEY2_GET1 =>
		SOURCE_REG <= SEL_IO;
		DEST_REG <= SEL_DES_LOW;
		NEWSTATE <= S_DES_KEY2_WAIT;
	    when S_DES_KEY2_WAIT =>
		if DATA_VALID = '0' then
		    NEWSTATE <= S_DES_KEY2_WAIT;
		else
		    NEWSTATE <= S_DES_KEY2_GET2;
		end if;
	    when S_DES_KEY2_GET2 =>
		SOURCE_REG <= SEL_IO;
		DEST_REG <= SEL_DES_HIGH;
		NEWSTATE <= S_DES_KEY2_WRITE;
	    when S_DES_KEY2_WRITE =>
		DES_DATA_IS_KEY_I <= '1';
		DES_DATA_READY_SET <= '1';
		NEWSTATE <= S_DES_KEY2_WAIT2;
	    when S_DES_KEY2_WAIT2 => 
		if DES_DATA_READY = '1' then
		    NEWSTATE <= S_DES_KEY2_WAIT2;
		else
		    if CTRL(1 downto 0) /= "01" then
			NEWSTATE <= S_DES_KEY3;
		    else
			NEWSTATE <= S_DES_READ_WRITE;
		    end if;
		end if;
	    when S_DES_KEY3 =>
		if DES_DATA_READY = '1' or DATA_VALID = '0' then
		    NEWSTATE <= S_DES_KEY3;
		else
		    NEWSTATE <= S_DES_KEY3_GET1;
		end if;
	    when S_DES_KEY3_GET1 =>
		SOURCE_REG <= SEL_IO;
		DEST_REG <= SEL_DES_LOW;
		NEWSTATE <= S_DES_KEY3_WAIT;
	    when S_DES_KEY3_WAIT =>
		if DATA_VALID = '0' then
		    NEWSTATE <= S_DES_KEY3_WAIT;
		else
		    NEWSTATE <= S_DES_KEY3_GET2;
		end if;
	    when S_DES_KEY3_GET2 =>
		SOURCE_REG <= SEL_IO;
		DEST_REG <= SEL_DES_HIGH;
		NEWSTATE <= S_DES_KEY3_WRITE;
	    when S_DES_KEY3_WRITE =>
		DES_DATA_IS_KEY_I <= '1';
		DES_DATA_READY_SET <= '1';
		NEWSTATE <= S_DES_KEY3_WAIT2;
	    when S_DES_KEY3_WAIT2 => 
		if DES_DATA_READY = '1' then
		    NEWSTATE <= S_DES_KEY3_WAIT2;
		else
		    NEWSTATE <= S_DES_READ_WRITE;
		end if;
		
	    when S_DES_READ_WRITE =>
		DES_DATA_IS_KEY_I <= '0';
		if DES_DATA_READY = '0' and DATA_VALID = '1' then
		    NEWSTATE <= S_DES_WRITE_REG1;
		elsif DES_BUFFER_FREE='0' and DOUT_EMPTY = '1' then
		    NEWSTATE <= S_DES_READ_REG1;
		else
		    NEWSTATE <= S_DES_READ_WRITE;
		end if;
		
	    when S_DES_WRITE_REG1 =>
		SOURCE_REG <= SEL_IO;
		DEST_REG <= SEL_DES_LOW;
		NEWSTATE <= S_DES_WRITE_WAIT;
	    when S_DES_WRITE_WAIT =>
		if DATA_VALID = '0' then
		    NEWSTATE <= S_DES_WRITE_WAIT;		    
		else
		    NEWSTATE <= S_DES_WRITE_REG2;
		end if;
	    when S_DES_WRITE_REG2 =>
		SOURCE_REG <= SEL_IO;
		DEST_REG <= SEL_DES_HIGH;
		NEWSTATE <= S_DES_WRITE;
	    when S_DES_WRITE =>
		DES_DATA_READY_SET <= '1';
		NEWSTATE <= S_DES_READ_WRITE;

	    when S_DES_READ_REG1 =>
		SOURCE_REG <= SEL_DES_LOW;
		DEST_REG <= SEL_IO;
		NEWSTATE <= S_DES_READ_WAIT;
	    when S_DES_READ_WAIT =>
		if DOUT_EMPTY = '0' then
		    NEWSTATE <= S_DES_READ_WAIT;		    
		else
		    NEWSTATE <= S_DES_READ_REG2;
		end if;
	    when S_DES_READ_REG2 =>
		SOURCE_REG <= SEL_DES_HIGH;
		DEST_REG <= SEL_IO;
		NEWSTATE <= S_DES_READ;
	    when S_DES_READ =>
		DES_BUFFER_FREE_SET <= '1';
		NEWSTATE <= S_DES_READ_WRITE;

	    when S_AUTHENTIFY =>  	--  --  --  --  --
		DES_DATA_IS_KEY_I <= '1';
		NEWSTATE <= S_AUTHENTIFY_WAIT;
	    when S_AUTHENTIFY_WAIT =>
		if DATA_VALID = '1' then
		  if DES_DATA_READY = '0' then
		      NEWSTATE <= S_MAKE_SIG_WRITE1;
		  else
		      NEWSTATE <= S_MAKE_SIG_WAIT1B;
		  end if;		    
		else
		    NEWSTATE <= S_AUTHENTIFY_WAIT;
		end if;
		
	    when S_MAKE_SIGNAUTURE =>  	--  --  --  --  --
		SOURCE_REG <= SEL_LFSR_CONST;  -- dummy egal
		DEST_REG <= SEL_IO;  	-- flush output-buffer
		DES_DATA_IS_KEY_I <= '1';
		NEWSTATE <= S_MAKE_SIG_WAIT1A;
	    when S_MAKE_SIG_WAIT1A =>
		if DATA_VALID = '1' then
		  if DES_DATA_READY = '0' then
		      NEWSTATE <= S_MAKE_SIG_WRITE1A;
		  else
		      NEWSTATE <= S_MAKE_SIG_WAIT1B;
		  end if;		    
		elsif DOUT_EMPTY = '1' then
		    NEWSTATE <= S_MAKE_SIG_RSA_WAIT1;
		else
		    NEWSTATE <= S_MAKE_SIG_WAIT1A;
		end if;
	    when S_MAKE_SIG_WAIT1 =>
		if DATA_VALID = '1' then
		  if DES_DATA_READY = '0' then
		      NEWSTATE <= S_MAKE_SIG_WRITE1;
		  else
		      NEWSTATE <= S_MAKE_SIG_WAIT1B;
		  end if;		    
		elsif DOUT_EMPTY = '1' then
		    NEWSTATE <= S_MAKE_SIG_RSA_WAIT1;
		else
		    NEWSTATE <= S_MAKE_SIG_WAIT1;
		end if;
	    when S_MAKE_SIG_WAIT1B =>
		if DES_DATA_READY = '0' then
		    NEWSTATE <= S_MAKE_SIG_WRITE1;
		else
		    NEWSTATE <= S_MAKE_SIG_WAIT1B;
		end if;
	    when S_MAKE_SIG_WRITE1A =>
		SOURCE_REG <= SEL_IO;
		DEST_REG <= SEL_DES_LOW;
		NEWSTATE <= S_MAKE_SIG_WAIT2;
	    when S_MAKE_SIG_WRITE1 =>
		DES_DATA_IS_KEY_I <= '0';
		SOURCE_REG <= SEL_IO;
		DEST_REG <= SEL_DES_LOW;
		NEWSTATE <= S_MAKE_SIG_WAIT2;
	    when S_MAKE_SIG_WAIT2 =>
		if DATA_VALID = '0' then
		    NEWSTATE <= S_MAKE_SIG_WAIT2;
		else
		    NEWSTATE <= S_MAKE_SIG_WRITE2;
		end if;
	    when S_MAKE_SIG_WRITE2 =>
		RAM_MODE <= RAM_MODE_SET_TEMPEXP;
		DES_BUFFER_FREE_SET <= '1';
		SOURCE_REG <= SEL_IO;
		DEST_REG <= SEL_DES_HIGH;
		NEWSTATE <= S_MAKE_SIG_WRITE;
	    when S_MAKE_SIG_WRITE =>
		RAM_MODE <= RAM_MODE_INC;
		DES_DATA_READY_SET <= '1';
		if CTRL(4 downto 0) = "01011" then  -- signate
		    NEWSTATE <= S_MAKE_SIG_WAIT1;
		else
		    NEWSTATE <= S_MAKE_SIG_RSA_WAIT1;
		end if;
	    when S_MAKE_SIG_RSA_WAIT1 =>
		RSA_SEL_I <= RSA_SEL_DATA;
		if DES_BUFFER_FREE='0' then
		    if DES_DATA_READY = '0' then
			NEWSTATE <= S_MAKE_SIG_RSA_COPY1;
		    else
			NEWSTATE <= S_MAKE_SIG_RSA_IGNORE;
		    end if;
		else
		    NEWSTATE <= S_MAKE_SIG_RSA_WAIT1;
		end if;
	    when S_MAKE_SIG_RSA_IGNORE =>
		DES_BUFFER_FREE_SET <= '1';
		NEWSTATE <= S_MAKE_SIG_RSA_WAIT1;
	    when S_MAKE_SIG_RSA_COPY1 =>
		RAM_MODE <= RAM_MODE_INC;
		SOURCE_REG <= SEL_DES_LOW;
		DEST_REG <= SEL_RSA;
		NEWSTATE <= S_MAKE_SIG_RSA_WRITE1;
	    when S_MAKE_SIG_RSA_WRITE1 => 
		RSA_VAL_ACC <= '1';
		NEWSTATE <= S_MAKE_SIG_RSA_WAIT2;
	    when S_MAKE_SIG_RSA_WAIT2 => 
		if RSA_READY = '1' then
		    NEWSTATE <= S_MAKE_SIG_RSA_COPY2;
		else
		    NEWSTATE <= S_MAKE_SIG_RSA_WAIT2;
		end if;
	    when S_MAKE_SIG_RSA_COPY2 =>
		RAM_MODE <= RAM_MODE_INC;
		SOURCE_REG <= SEL_DES_HIGH;
		DEST_REG <= SEL_RSA;
		NEWSTATE <= S_MAKE_SIG_RSA_WRITE2;
	    when S_MAKE_SIG_RSA_WRITE2 => 
		RSA_VAL_ACC <= '1';
		NEWSTATE <= S_MAKE_SIG_RSA_WAIT3;
	    when S_MAKE_SIG_RSA_WAIT3 => 
		if RSA_READY = '1' then
		    NEWSTATE <= S_MAKE_SIG_RSA_LFSR_COPY;
		else
		    NEWSTATE <= S_MAKE_SIG_RSA_WAIT3;
		end if;
	    when S_MAKE_SIG_RSA_LFSR_COPY =>
		RAM_MODE <= RAM_MODE_INC;
		SOURCE_REG <= SEL_LFSR_LOW;
		DEST_REG <= SEL_RSA;
		NEWSTATE <= S_MAKE_SIG_RSA_LFSR_WRITE;
	    when S_MAKE_SIG_RSA_LFSR_WRITE => 
		RSA_VAL_ACC <= '1';
		NEWSTATE <= S_MAKE_SIG_RSA_LFSR_WAIT;
	    when S_MAKE_SIG_RSA_LFSR_WAIT => 
		if RSA_READY = '1' then
		    if RAM_ADR_IS_AT_END_OFF_TEMPEXP /= '1' then
			NEWSTATE <= S_MAKE_SIG_RSA_LFSR_COPY;
		    else
			NEWSTATE <= S_MAKE_SIG_RSA_COPY4;
		    end if;
		else
		    NEWSTATE <= S_MAKE_SIG_RSA_LFSR_WAIT;
		end if;
	    when S_MAKE_SIG_RSA_COPY4 =>
		SOURCE_REG <= SEL_LFSR_CONST;
		DEST_REG <= SEL_RSA;
		RSA_VAL_ACC <= '1';
		NEWSTATE <= S_DECRYPT_RSA;

	    when S_CHECK_SIGNATURE =>  	--  --  --  --  --
		RESULT_I <= '0';
		NEWSTATE <= S_ENCRYPT_RSA;  ---> RSA
	    when S_CHECKSIGN_RSAREAD =>
		SOURCE_REG <= SEL_LFSR_LOW;  -- set out buffer full
		DEST_REG <= SEL_IO;
		RSA_SEL_I <= RSA_SEL_READ;
		RAM_MODE <= RAM_MODE_SET_DES_KEY;
		if RSA_READY='1' then
		    NEWSTATE <= S_CHECKSIGN_RSAREAD_COPY1;
		else
		    NEWSTATE <= S_CHECKSIGN_RSAREAD;
		end if;
	    when S_CHECKSIGN_RSAREAD_COPY1 =>
		RAM_MODE <= RAM_MODE_INC;
		SOURCE_REG <= SEL_RSA;
		DEST_REG <= SEL_RAM;
		RSA_VAL_ACC <= '1';
		NEWSTATE <= S_CHECKSIGN_RSAREAD_WAIT2;
	    when S_CHECKSIGN_RSAREAD_WAIT2 =>
		if RSA_READY = '1' then
		    NEWSTATE <= S_CHECKSIGN_RSAREAD_COPY2;
		else
		    NEWSTATE <= S_CHECKSIGN_RSAREAD_WAIT2;
		end if;
	    when S_CHECKSIGN_RSAREAD_COPY2 =>
		SOURCE_REG <= SEL_RSA;
		DEST_REG <= SEL_RAM;
		RSA_VAL_ACC <= '1';
		DES_DATA_IS_KEY_I <= '1';
		NEWSTATE <= S_CHECKSIGN_HASH;
	    when S_CHECKSIGN_HASH =>
		if DOUT_EMPTY = '1' then
		    NEWSTATE <= S_CHECKSIGN_ISEQ_LOW_LOAD;
		elsif DATA_VALID = '1' then
		  if DES_DATA_READY = '0' then
		      NEWSTATE <= S_CHECKSIGN_HASH_WRITE1;
		  else
		      NEWSTATE <= S_CHECKSIGN_HASH_WAIT1B;
		  end if;
		else
		    NEWSTATE <= S_CHECKSIGN_HASH;
		end if;
	    when S_CHECKSIGN_HASH_WAIT1B =>
		RESULT_I <= '0';
		if DES_DATA_READY = '0' then
		    NEWSTATE <= S_CHECKSIGN_HASH_WRITE1;
		else
		    NEWSTATE <= S_CHECKSIGN_HASH_WAIT1B;
		end if;
	    when S_CHECKSIGN_HASH_WRITE1 =>
		RESULT_I <= '0';
		SOURCE_REG <= SEL_IO;
		DEST_REG <= SEL_DES_LOW;
		NEWSTATE <= S_CHECKSIGN_HASH_WAIT2;
	    when S_CHECKSIGN_HASH_WAIT2 =>
		if DATA_VALID = '0' then
		    NEWSTATE <= S_CHECKSIGN_HASH_WAIT2;
		else
		    NEWSTATE <= S_CHECKSIGN_HASH_WRITE2;
		end if;
	    when S_CHECKSIGN_HASH_WRITE2 =>
		DES_BUFFER_FREE_SET <= '1';
		SOURCE_REG <= SEL_IO;
		DEST_REG <= SEL_DES_HIGH;
		NEWSTATE <= S_CHECKSIGN_HASH_WRITE;
	    when S_CHECKSIGN_HASH_WRITE =>
		DES_DATA_READY_SET <= '1';
		NEWSTATE <= S_CHECKSIGN_HASH_WAIT3;
	    when S_CHECKSIGN_HASH_WAIT3 =>
		RAM_MODE <= RAM_MODE_SET_DES_KEY;
		if DES_BUFFER_FREE='0' then
		    NEWSTATE <= S_CHECKSIGN_HASH_NOKEY;
		else
		    NEWSTATE <= S_CHECKSIGN_HASH_WAIT3;
		end if;
	    when S_CHECKSIGN_HASH_NOKEY =>
		DES_DATA_IS_KEY_I <= '0';
		NEWSTATE <= S_CHECKSIGN_HASH;
	    when S_CHECKSIGN_ISEQ_LOW_LOAD =>
		DES_DATA_IS_KEY_I <= '0';
		SOURCE_REG <= SEL_RAM;  --1
		NEWSTATE <= S_CHECKSIGN_ISEQ_LOW_CHECK_RAMACCESS;
	    when S_CHECKSIGN_ISEQ_LOW_CHECK_RAMACCESS =>
		RAM_MODE <= RAM_MODE_INC;
		SOURCE_REG <= SEL_RAM;  --2
		EQ_REG <= '1';
		NEWSTATE <= S_CHECKSIGN_ISEQ_LOW_CHECK;
	    when S_CHECKSIGN_ISEQ_LOW_CHECK =>
		SOURCE_REG <= SEL_DES_LOW;
		NEWSTATE <= S_CHECKSIGN_ISEQ_LOW_JUMP;
	    when S_CHECKSIGN_ISEQ_LOW_JUMP =>
		if EQUAL = '1' then
		    NEWSTATE <= S_CHECKSIGN_ISEQ_HIGH_LOAD;
		else
		    NEWSTATE <= S_IDLE;
		end if;
	    when S_CHECKSIGN_ISEQ_HIGH_LOAD =>
		SOURCE_REG <= SEL_RAM;  --1
		EQ_REG <= '1';
		NEWSTATE <= S_CHECKSIGN_ISEQ_HIGH_CHECK_RAMACCESS;
	    when S_CHECKSIGN_ISEQ_HIGH_CHECK_RAMACCESS =>
		SOURCE_REG <= SEL_RAM;  --2
		EQ_REG <= '1';
		NEWSTATE <= S_CHECKSIGN_ISEQ_HIGH_CHECK;
	    when S_CHECKSIGN_ISEQ_HIGH_CHECK =>
		SOURCE_REG <= SEL_DES_HIGH;
		NEWSTATE <= S_CHECKSIGN_ISEQ_HIGH_JUMP;
	    when S_CHECKSIGN_ISEQ_HIGH_JUMP =>
		if EQUAL = '1' then
		    NEWSTATE <= S_CHECKSIGN_ISEQ_OK;
		else
		    NEWSTATE <= S_IDLE;
		end if;
	    when S_CHECKSIGN_ISEQ_OK =>
		RESULT_I <= '1';
		NEWSTATE <= S_IDLE;

		
	    when S_CHECK_AUTHENTIFY =>  --  --  --  --  --
		RESULT_I <= '0';  	      -- get a random key
		RAM_MODE <= RAM_MODE_SET_DES_KEY;
		NEWSTATE <= S_CHECKAUTH_PREHASH_WAIT;
	    when S_CHECKAUTH_PREHASH_WAIT =>  -- make in nearly random with DES
		if DES_DATA_READY='0' then
		    NEWSTATE <= S_CHECKAUTH_PREHASH_COPY_L;
		else
		    NEWSTATE <= S_CHECKAUTH_PREHASH_WAIT;
		end if;
	    when S_CHECKAUTH_PREHASH_COPY_L =>
		SOURCE_REG <= SEL_LFSR_LOW;
		DEST_REG <= SEL_DES_LOW;
		NEWSTATE <= S_CHECKAUTH_PREHASH_COPY_H;
	    when S_CHECKAUTH_PREHASH_COPY_H =>
		SOURCE_REG <= SEL_LFSR_HIGH;
		DEST_REG <= SEL_DES_HIGH;
		DES_DATA_READY_SET <= '1';
		DES_DATA_IS_KEY_I <= '1';
		NEWSTATE <= S_CHECKAUTH_PREHASH_WAIT2;
	    when S_CHECKAUTH_PREHASH_WAIT2 =>
		if DES_BUFFER_FREE='0' then
		    NEWSTATE <= S_CHECKAUTH_PREHASH_COPYBACK_L;
		else
		    NEWSTATE <= S_CHECKAUTH_PREHASH_WAIT2;
		end if;
	    when S_CHECKAUTH_PREHASH_COPYBACK_L =>
		RAM_MODE <= RAM_MODE_INC;
		SOURCE_REG <= SEL_DES_LOW;
		DEST_REG <= SEL_RAM;
		NEWSTATE <= S_CHECKAUTH_PREHASH_COPYBACK_H;
	    when S_CHECKAUTH_PREHASH_COPYBACK_H =>
		RAM_MODE <= RAM_MODE_SET_DES_KEY;
		SOURCE_REG <= SEL_DES_HIGH;
		DEST_REG <= SEL_RAM;
		DES_BUFFER_FREE_SET <= '1';
		NEWSTATE <= S_CHECKAUTH_OL_WAIT;
	    when S_CHECKAUTH_OL_WAIT =>  -- send random key to other
		if DOUT_EMPTY='1' then
		    NEWSTATE <= S_CHECKAUTH_OL_COPY;
		else
		    NEWSTATE <= S_CHECKAUTH_OL_WAIT;
		end if;
	    when S_CHECKAUTH_OL_COPY =>
		SOURCE_REG <= SEL_RAM; --1
		NEWSTATE <= S_CHECKAUTH_OH_WAIT_RAMACCESS;
	    when S_CHECKAUTH_OH_WAIT_RAMACCESS =>
		RAM_MODE <= RAM_MODE_INC;
		SOURCE_REG <= SEL_RAM; --2
		DEST_REG <= SEL_IO;
		NEWSTATE <= S_CHECKAUTH_OH_WAIT;
	    when S_CHECKAUTH_OH_WAIT =>
		if DOUT_EMPTY='1' then
		    NEWSTATE <= S_CHECKAUTH_OH_COPY;
		else
		    NEWSTATE <= S_CHECKAUTH_OH_WAIT;
		end if;
	    when S_CHECKAUTH_OH_COPY =>
		SOURCE_REG <= SEL_RAM; --1
		NEWSTATE <= S_CHECKAUTH_HASH_WAIT_RAMACCESS;
	    when S_CHECKAUTH_HASH_WAIT_RAMACCESS =>
		RAM_MODE <= RAM_MODE_SET_DES_KEY;
		SOURCE_REG <= SEL_RAM; --2
		DEST_REG <= SEL_IO;
		NEWSTATE <= S_CHECKAUTH_HASH_WAIT;
	    when S_CHECKAUTH_HASH_WAIT =>  -- put random key into des
		if DES_DATA_READY='0' then
		    NEWSTATE <= S_CHECKAUTH_HASH_COPY_L;
		else
		    NEWSTATE <= S_CHECKAUTH_HASH_WAIT;
		end if;
	    when S_CHECKAUTH_HASH_COPY_L =>
		SOURCE_REG <= SEL_RAM; --1
		NEWSTATE <= S_CHECKAUTH_HASH_COPY_H_RAMACCESS;
	    when S_CHECKAUTH_HASH_COPY_H_RAMACCESS =>
		RAM_MODE <= RAM_MODE_INC;
		SOURCE_REG <= SEL_RAM; --2
		DEST_REG <= SEL_DES_LOW;
		NEWSTATE <= S_CHECKAUTH_HASH_COPY_H;
	    when S_CHECKAUTH_HASH_COPY_H =>
		SOURCE_REG <= SEL_RAM;  --1
		NEWSTATE <= S_CHECKAUTH_HASH_WAIT2_RAMACCESS;
	    when S_CHECKAUTH_HASH_WAIT2_RAMACCESS =>
		RAM_MODE <= RAM_MODE_SET_DES_KEY;
		SOURCE_REG <= SEL_RAM;  --2
		DEST_REG <= SEL_DES_HIGH;
		DES_DATA_IS_KEY_I <= '1';
		DES_DATA_READY_SET <= '1';
		NEWSTATE <= S_CHECKAUTH_HASH_WAIT2;
	    when S_CHECKAUTH_HASH_WAIT2 =>
		if DES_BUFFER_FREE='0' then
		    NEWSTATE <= S_CHECKAUTH_HASH_COPYBACK_L;
		else
		    NEWSTATE <= S_CHECKAUTH_HASH_WAIT2;
		end if;
	    when S_CHECKAUTH_HASH_COPYBACK_L =>
		RAM_MODE <= RAM_MODE_INC;
		SOURCE_REG <= SEL_DES_LOW;
		DEST_REG <= SEL_RAM;
		NEWSTATE <= S_CHECKAUTH_HASH_COPYBACK_H;
	    when S_CHECKAUTH_HASH_COPYBACK_H =>
		SOURCE_REG <= SEL_DES_HIGH;
		DEST_REG <= SEL_RAM;
		NEWSTATE <= S_ENCRYPT_RSA; ---> RSA
	    when S_CHECKAUTH_RRSA_WAIT1 =>  -- compare encrypted with DES result
		RSA_SEL_I <= RSA_SEL_READ;
		RAM_MODE <= RAM_MODE_SET_DES_KEY;
		if RSA_READY = '1' then
		    NEWSTATE <= S_CHECKAUTH_RRSA_WORD1;
		else
		    NEWSTATE <= S_CHECKAUTH_RRSA_WAIT1;
		end if;
	    when S_CHECKAUTH_RRSA_WORD1 =>
		SOURCE_REG <= SEL_RSA;
		EQ_REG  <= '1';
		NEWSTATE <= S_CHECKAUTH_RRSA_CHECK;
	    when S_CHECKAUTH_RRSA_CHECK =>
		SOURCE_REG <= SEL_RAM;  --1
		NEWSTATE <= S_CHECKAUTH_RRSA_CHECK_RAMACCESS;
	    when S_CHECKAUTH_RRSA_CHECK_RAMACCESS =>
		RAM_MODE <= RAM_MODE_INC;
		SOURCE_REG <= SEL_RAM;  --2
		NEWSTATE <= S_CHECKAUTH_RRSA_WAIT2;
	    when S_CHECKAUTH_RRSA_WAIT2 =>
	        RSA_VAL_ACC <= '1';
		if EQUAL = '1' then
		    if RSA_READY = '0' then
			NEWSTATE <= S_CHECKAUTH_RRSA_WAIT2B;
		    else
			NEWSTATE <= S_CHECKAUTH_RRSA_WORD2;
		    end if;
		else
		    NEWSTATE <= S_IDLE;
		end if;
	    when S_CHECKAUTH_RRSA_WAIT2B =>
		if RSA_READY = '0' then
		    NEWSTATE <= S_CHECKAUTH_RRSA_WAIT2B;
		else
		    NEWSTATE <= S_CHECKAUTH_RRSA_WORD2;
		end if;
	    when S_CHECKAUTH_RRSA_WORD2 =>
	        RSA_VAL_ACC <= '1';
		SOURCE_REG <= SEL_RSA;
		EQ_REG <= '1';
		NEWSTATE <= S_CHECKAUTH_RRSA_DECIDE;
	    when S_CHECKAUTH_RRSA_DECIDE =>
		SOURCE_REG <= SEL_RAM;  --1
		NEWSTATE <= S_CHECKAUTH_RRSA_DECIDE_RAMACCESS;
	    when S_CHECKAUTH_RRSA_DECIDE_RAMACCESS =>
		SOURCE_REG <= SEL_RAM;  --2
		NEWSTATE <= S_CHECKAUTH_RRSA_JUMP;
	    when S_CHECKAUTH_RRSA_JUMP =>
		if EQUAL = '1' then
		    if RESULT_I = '1' then
			NEWSTATE <= S_CHECKAUTH_OK2;
		    else
			NEWSTATE <= S_CHECKAUTH_OK;
		    end if;
		else
		    NEWSTATE <= S_IDLE;
		end if;
	    when S_CHECKAUTH_OK =>  	-- Yes it is EQ
		RESULT_I <= '1';
		RAM_MODE <= RAM_MODE_SET_TEMPEXP;
		if DES_DATA_READY='0' then
		    NEWSTATE <= S_CHECKAUTH_HASH2_COPY_L;
		else
		    NEWSTATE <= S_CHECKAUTH_OK;
		end if;
	    when S_CHECKAUTH_HASH2_COPY_L =>  -- DES-hash over first 64bit of RSA-key
		SOURCE_REG <= SEL_RAM;  --1
		NEWSTATE <= S_CHECKAUTH_HASH2_COPY_L_RAMACCESS;
	    when S_CHECKAUTH_HASH2_COPY_L_RAMACCESS =>
		RAM_MODE <= RAM_MODE_INC;
		SOURCE_REG <= SEL_RAM;  --2
		DEST_REG <= SEL_DES_LOW;
		NEWSTATE <= S_CHECKAUTH_HASH2_COPY_H;
	    when S_CHECKAUTH_HASH2_COPY_H =>
		SOURCE_REG <= SEL_RAM;  --1
		NEWSTATE <= S_CHECKAUTH_HASH2_COPY_H_RAMACCESS;
	    when S_CHECKAUTH_HASH2_COPY_H_RAMACCESS =>
		RAM_MODE <= RAM_MODE_INC;
		SOURCE_REG <= SEL_RAM;  --2
		DEST_REG <= SEL_DES_HIGH;
		DES_DATA_READY_SET <= '1';
		DES_DATA_IS_KEY_I <= '1';  -- first is a key
		DES_BUFFER_FREE_SET <= '1';
		NEWSTATE <= S_CHECKAUTH_HASH2_WAIT;
	    when S_CHECKAUTH_HASH2_WAIT =>
		if DES_DATA_READY = '0' then
		    NEWSTATE <= S_CHECKAUTH_HASH2_COPY2_L;
		else
		    NEWSTATE <= S_CHECKAUTH_HASH2_WAIT;
		end if;
	    when S_CHECKAUTH_HASH2_COPY2_L =>  -- DES-hash over rest of RSA-key
		SOURCE_REG <= SEL_RAM;  --1
		NEWSTATE <= S_CHECKAUTH_HASH2_COPY2_L_RAMACCESS;
	    when S_CHECKAUTH_HASH2_COPY2_L_RAMACCESS =>
		RAM_MODE <= RAM_MODE_INC;
		SOURCE_REG <= SEL_RAM;  --2
		DEST_REG <= SEL_DES_LOW;
		NEWSTATE <= S_CHECKAUTH_HASH2_COPY2_H;
	    when S_CHECKAUTH_HASH2_COPY2_H =>
		SOURCE_REG <= SEL_RAM;  --1
		NEWSTATE <= S_CHECKAUTH_HASH2_COPY2_H_RAMACCESS;
	    when S_CHECKAUTH_HASH2_COPY2_H_RAMACCESS =>
		RAM_MODE <= RAM_MODE_INC;
		SOURCE_REG <= SEL_RAM;  --2
		DEST_REG <= SEL_DES_HIGH;
		DES_DATA_READY_SET <= '1';
		DES_DATA_IS_KEY_I <= '0';  -- rest is not a key
		DES_BUFFER_FREE_SET <= '1';
		NEWSTATE <= S_CHECKAUTH_HASH2_WAIT2;
	    when S_CHECKAUTH_HASH2_WAIT2 =>
		if (DES_DATA_READY = '0') AND (RAM_ADR_IS_AT_END_OFF_TEMPEXP /= '1') then
		    NEWSTATE <= S_CHECKAUTH_HASH2_COPY2_L;
		elsif (DES_BUFFER_FREE = '0') AND (RAM_ADR_IS_AT_END_OFF_TEMPEXP = '1' ) then
		    if DES_DATA_READY = '1' then
			NEWSTATE <= S_CHECKAUTH_HASH2_IGNORE;
		    else			
			NEWSTATE <= S_CHECKAUTH_HASH2_COPYBACK;			
		    end if;
		else
		    NEWSTATE <= S_CHECKAUTH_HASH2_WAIT2;
		end if;
	    when S_CHECKAUTH_HASH2_IGNORE =>
		DES_BUFFER_FREE_SET <= '1';
		NEWSTATE <= S_CHECKAUTH_HASH2_WAIT2;
	    when S_CHECKAUTH_HASH2_COPYBACK =>
		RAM_MODE <= RAM_MODE_SET_DES_KEY;
		NEWSTATE <= S_CHECKAUTH_HASH2_COPYBACK_L;
	    when S_CHECKAUTH_HASH2_COPYBACK_L =>
		RAM_MODE <= RAM_MODE_INC;
		SOURCE_REG <= SEL_DES_LOW;
		DEST_REG <= SEL_RAM;
		NEWSTATE <= S_CHECKAUTH_HASH2_COPYBACK_H;
	    when S_CHECKAUTH_HASH2_COPYBACK_H =>
		RSA_SEL_I <= RSA_SEL_MODULO;
		RAM_MODE <= RAM_MODE_SET_ZERTMODUL;
		SOURCE_REG <= SEL_DES_HIGH;
		DEST_REG <= SEL_RAM;
		DES_BUFFER_FREE_SET <= '1';
		NEWSTATE <= S_CHECKAUTH_RSA_MODUL_COPY;
	    when S_CHECKAUTH_RSA_MODUL_COPY => -- RSA with ZERT-key
		SOURCE_REG <= SEL_RAM;  --1
		NEWSTATE <= S_CHECKAUTH_RSA_MODUL_COPY_RAMACCESS;
	    when S_CHECKAUTH_RSA_MODUL_COPY_RAMACCESS =>
		RAM_MODE <= RAM_MODE_INC;
		SOURCE_REG <= SEL_RAM;  --2
		DEST_REG <= SEL_RSA;
		NEWSTATE <= S_CHECKAUTH_RSA_MODUL_WRITE;
	    when S_CHECKAUTH_RSA_MODUL_WRITE => 
		RSA_VAL_ACC <= '1';
		NEWSTATE <= S_CHECKAUTH_RSA_MODUL_WAIT;
	    when S_CHECKAUTH_RSA_MODUL_WAIT =>
		if RSA_READY = '0' then
		    NEWSTATE <= S_CHECKAUTH_RSA_MODUL_WAIT;
		else
		    if RAM_ADR_IS_AT_END_OFF_ZERTMODUL /= '1' then
			NEWSTATE <= S_CHECKAUTH_RSA_MODUL_COPY;
		    else
			NEWSTATE <= S_RSA_DATA_BEGIN; --------->
		    end if;
		end if;
	    when S_CHECKAUTH_OK2 =>
		SECURITY <= AUTHENTIFIED;
		NEWSTATE <= S_IDLE;
		
	    when S_SET_PIN  =>  	--  --  --  --  --
		RAM_MODE  <= RAM_MODE_SET_PIN;
      		if DATA_VALID='1' then
		    NEWSTATE <= S_SET_PIN_LOAD;
		else
		    NEWSTATE <= S_SET_PIN;
		end if;
	    when S_SET_PIN_LOAD =>
		SOURCE_REG <= SEL_IO;
		DEST_REG  <= SEL_RAM;
		NEWSTATE <= S_IDLE;


	    when S_SET_ZERT =>  	--  --  --  --  --
		RAM_MODE <= RAM_MODE_SET_ZERT;
		NEWSTATE <= S_SET_ZERT_WAIT;
	    when S_SET_ZERT_WAIT =>
		if DATA_VALID='1' then
		    NEWSTATE <= S_SET_ZERT_COPY;
		else
		    NEWSTATE <= S_SET_ZERT_WAIT;
		end if;
	    when S_SET_ZERT_COPY =>
		SOURCE_REG <= SEL_IO;
		DEST_REG <= SEL_RAM;
		RAM_MODE <= RAM_MODE_INC;
		NEWSTATE <= S_SET_ZERT_END;
	    when S_SET_ZERT_END =>
		if RAM_ADR_IS_AT_END_OFF_ZERTMODUL /= '1' then
		    NEWSTATE <= S_SET_ZERT_WAIT;
		else
		    NEWSTATE <= S_IDLE;
		end if;

		
	    when S_READ_PUBLIC_KEYS =>  --  --  --  --  --
		RAM_MODE <= RAM_MODE_SET_PUBLICKEY;
		NEWSTATE <= S_READ_PUBLIC_KEYS_WAIT;
	    when S_READ_PUBLIC_KEYS_WAIT =>
		if DOUT_EMPTY='1' then
		    NEWSTATE <= S_READ_PUBLIC_KEYS_COPY;
		else
		    NEWSTATE <= S_READ_PUBLIC_KEYS_WAIT;
		end if;
	    when S_READ_PUBLIC_KEYS_COPY =>
		SOURCE_REG <= SEL_RAM;  --1
		NEWSTATE <= S_READ_PUBLIC_KEYS_COPY_RAMACCESS;
	    when S_READ_PUBLIC_KEYS_COPY_RAMACCESS =>
		SOURCE_REG <= SEL_RAM;  --2
		DEST_REG <= SEL_IO;
		NEWSTATE <= S_READ_PUBLIC_KEYS_NEXT;
	    when S_READ_PUBLIC_KEYS_NEXT =>
		RAM_MODE <= RAM_MODE_INC;
		NEWSTATE <= S_READ_PUBLIC_KEYS_END;
	    when S_READ_PUBLIC_KEYS_END =>
		if RAM_ADR_IS_AT_END_OFF_PUBLICKEY = '1' then
		    NEWSTATE <= S_READ_PUBLIC_KEYS_NEXT2;		    
                elsif RAM_ADR_IS_AT_END_OFF_ZERTMODUL = '1' then
		    NEWSTATE <= S_IDLE;
		else
		    NEWSTATE <= S_READ_PUBLIC_KEYS_WAIT;
		end if;
	    when S_READ_PUBLIC_KEYS_NEXT2 =>
		RAM_MODE <= RAM_MODE_SET_MODUL;
		NEWSTATE <= S_READ_PUBLIC_KEYS_WAIT;
		
	    when S_READ_USER_DATA =>  	--  --  --  --  --
		RAM_MODE <= RAM_MODE_SET_USER;
		NEWSTATE <= S_READ_USER_DATA_WAIT;
	    when S_READ_USER_DATA_WAIT =>
		if DOUT_EMPTY='1' then
		    NEWSTATE <= S_READ_USER_DATA_COPY;
		else
		    NEWSTATE <= S_READ_USER_DATA_WAIT;
		end if;
	    when S_READ_USER_DATA_COPY =>
		SOURCE_REG <= SEL_RAM;  --1
		NEWSTATE <= S_READ_USER_DATA_COPY_RAMACCES;
	    when S_READ_USER_DATA_COPY_RAMACCES =>
		SOURCE_REG <= SEL_RAM;  --2
		DEST_REG <= SEL_IO;
		NEWSTATE <= S_READ_USER_DATA_NEXT;
	    when S_READ_USER_DATA_NEXT =>
		RAM_MODE <= RAM_MODE_INC;
		NEWSTATE <= S_READ_USER_DATA_END;
	    when S_READ_USER_DATA_END =>
		if RAM_ADR_IS_AT_END_OFF_ALL /= '1' then
		    NEWSTATE <= S_READ_USER_DATA_WAIT;
                else
		    NEWSTATE <= S_IDLE;
		end if;

	    when S_NAME_OUT =>
		RAM_SEL <= '1';
		RAM_MODE <= RAM_MODE_SET_PUBLICKEY;
		NEWSTATE <= S_NAME_OUT_COPY;
	    when S_NAME_OUT_COPY =>
		RAM_SEL <= '1';
		RAM_MODE <= RAM_MODE_INC;
		SOURCE_REG <= SEL_RAM;	-- NAME ROM
		DEST_REG <= SEL_IO;
		NEWSTATE <= S_NAME_OUT_NEXT;
	    when S_NAME_OUT_NEXT =>
		RAM_SEL <= '1';
		if DOUT_EMPTY = '0' then
		    NEWSTATE <= S_NAME_OUT_NEXT;
		else
		    NEWSTATE <= S_NAME_OUT_COPY;
		end if;

	    when S_RAMTEST_WAIT_EXPECTED =>
	        RESULT_I <= '1';
		RAM_MODE <= RAM_MODE_SET_PUBLICKEY;
		if DATA_VALID = '1' then
		    NEWSTATE <= S_RAMTEST_COPY_EXPECTED;
		else
		    NEWSTATE <= S_RAMTEST_WAIT_EXPECTED;
		end if;
	    when S_RAMTEST_COPY_EXPECTED =>
		SOURCE_REG <= SEL_IO;
		EQ_REG <= '1';
		NEWSTATE <= S_RAMTEST_WAIT_DATA;
	    when S_RAMTEST_WAIT_DATA =>
		SOURCE_REG <= SEL_RAM;  --1
		if DATA_VALID = '1' then
		    NEWSTATE <= S_RAMTEST_CHECK;
		else
		    NEWSTATE <= S_RAMTEST_WAIT_DATA;
		end if;
	    when S_RAMTEST_CHECK =>
		SOURCE_REG <= SEL_RAM;  --2
		NEWSTATE <= S_RAMTEST_WRITE;
	    when S_RAMTEST_WRITE =>
		RAM_MODE <= RAM_MODE_INC;
		SOURCE_REG <= SEL_IO;
		DEST_REG <= SEL_RAM;
		if EQUAL = '0' then
		    NEWSTATE <= S_RAMTEST_FAIL;
		else
		    NEWSTATE <= S_RAMTEST_NEXT;
		end if;
	    when S_RAMTEST_FAIL =>
		RESULT_I <= '0';
		NEWSTATE <= S_RAMTEST_NEXT;
	    when S_RAMTEST_NEXT =>
		SOURCE_REG <= SEL_RAM;  --1
		if RAM_ADR_IS_AT_END_OFF_ALL = '1' then
		    NEWSTATE <= S_IDLE;
		else
		    NEWSTATE <= S_RAMTEST_CHECK;
		end if;
		
            -- idle --
            when S_IDLE =>
		NEWSTATE <= S_IDLE;
		
	    -- others --
	    when others =>
		NEWSTATE <= S_RESET;
	end case;
    end process;

    DES_DATA_IS_KEY <= DES_DATA_IS_KEY_I;
    RSA_SEL <= RSA_SEL_I;
    
    DES_IN_EN <= DES_BUFFER_FREE;
    DES_MODE(4 downto 0) <= CTRL(4 downto 0);

    INVERT <= CTRL(6) when SECURITY=NO_KEY else '0';

    INT <= ( not DOUT_EMPTY ) and CTRL(7);

    ENABLE_TEST <=  not ( SECURITY(0) or SECURITY(1) );

    STATUS(7) <= '1' when STATE=S_IDLE else '0';  -- nothing to do
    STATUS(6) <= '1' when STATE<S_NEWCOMMAND else '0';  -- insecure
    STATUS(5) <= DES_ERR;  			-- TEST ??
    STATUS(4) <= DES_PARITY;  		-- DES?-Key-Paryty? ERROR
    STATUS(3) <= '1' when SECURITY=AUTHENTIFIED else '0';
    STATUS(2) <= RESULT_I;		-- The result of a check-command.
    STATUS(1) <= not DOUT_EMPTY;  	-- Data-out buffer is full. (user can read)
    STATUS(0) <= not DATA_VALID;  	-- Data-in  buffer is empty. (user can write)
    
end BEHAVIORAL;


library IEEE;
   use IEEE.std_logic_1164.all;
   use IEEE.std_logic_misc.all;
   use WORK.RAM_ADR_CONST.all;

entity FSM is
      Port ( CARDCHANGE : In    std_logic;
	     CLK : In    std_logic;
	     CTRL : In    std_logic_vector (7 downto 0);
             CTRL_CHANGE : In    std_logic;
             DATA_VALID : In    std_logic;
             DES_BUFFER_FREE : In    std_logic;
             DES_DATA_READY : In    std_logic;
             DES_ERR : In    std_logic;
             DES_PARITY : In    std_logic;
             DOUT_EMPTY : In    std_logic;
	     EQUAL : In    std_logic;
	     RESET : In    std_logic;
             RSA_NEXTEXP : In    std_logic;
             RSA_READY : In    std_logic;
             BUSY : Out   std_logic;
             DES_BUFFER_FREE_SET : Out   std_logic;
             DES_DATA_IS_KEY : Out   std_logic;
             DES_DATA_READY_SET : Out   std_logic;
             DES_IN_EN : Out   std_logic;
             DES_MODE : Out   std_logic_vector (4 downto 0);
             DEST_REG : Out   std_logic_vector (2 downto 0);
             ENABLE_TEST : Out   std_logic;
             EQ_REG : Out   std_logic;
             INT : Out   std_logic;
             RAM_ADR : Out   std_logic_vector (7 downto 0);
             RAM_SEL : Out   std_logic;
             RSA_GO : Out   std_logic;
             RSA_SEL : Out   std_logic_vector (1 downto 0);
             RSA_VAL_ACC : Out   std_logic;
             SOURCE_REG : Out   std_logic_vector (2 downto 0);
             STATE_EN : Out   std_logic;
             STATUS : Out   std_logic_vector (7 downto 0) );
end FSM;

architecture BEHAVIORAL of FSM is

    component RAM_COUNTER
	port ( RAM_ADR : out STD_LOGIC_VECTOR(7 downto 0);
	       CLK : in STD_LOGIC;  	-- clock
	       RESET : in STD_LOGIC;  	-- reset
	       RAM_MODE : in STD_LOGIC_VECTOR(5 downto 0);
	       RAM_ADR_IS_AT_END_OFF_ALL		: Out   std_logic;
	       RAM_ADR_IS_AT_END_OFF_TEMPEXP	: Out   std_logic;
	       RAM_ADR_IS_AT_END_OFF_MODUL		: Out   std_logic;
	       RAM_ADR_IS_AT_END_OFF_PUBLICKEY	: Out   std_logic;
	       RAM_ADR_IS_AT_END_OFF_PRIVATKEY	: Out   std_logic;
	       RAM_ADR_IS_AT_END_OFF_ZERTPUB	: Out   std_logic;
	       RAM_ADR_IS_AT_END_OFF_ZERTMODUL	: Out   std_logic;
	       INVERT : in STD_LOGIC );
    end component;

    component FSM_CORE
      Port ( CARDCHANGE : In    std_logic;
	     CLK : In    std_logic;
	     CTRL : In    std_logic_vector (7 downto 0);
             CTRL_CHANGE : In    std_logic;
             DATA_VALID : In    std_logic;
             DES_BUFFER_FREE : In    std_logic;
             DES_DATA_READY : In    std_logic;
             DES_ERR : In    std_logic;
             DES_PARITY : In    std_logic;
             DOUT_EMPTY : In    std_logic;
	     EQUAL : In    std_logic;
	     RESET : In    std_logic;
             RSA_NEXTEXP : In    std_logic;
             RSA_READY : In    std_logic;
             BUSY : Out   std_logic;
             DES_BUFFER_FREE_SET : Out   std_logic;
             DES_DATA_IS_KEY : Out   std_logic;
             DES_DATA_READY_SET : Out   std_logic;
             DES_IN_EN : Out   std_logic;
             DES_MODE : Out   std_logic_vector (4 downto 0);
             DEST_REG : Out   std_logic_vector (2 downto 0);
             ENABLE_TEST : Out   std_logic;
             EQ_REG : Out   std_logic;
             INT : Out   std_logic;
             RAM_SEL : Out   std_logic;
             RSA_GO : Out   std_logic;
             RSA_SEL : Out   std_logic_vector (1 downto 0);
             RSA_VAL_ACC : Out   std_logic;
             SOURCE_REG : Out   std_logic_vector (2 downto 0);
             STATE_EN : Out   std_logic;
             STATUS : Out   std_logic_vector (7 downto 0);
	     RAM_MODE : Out STD_LOGIC_VECTOR(5 downto 0);
	     RAM_ADR_IS_AT_END_OFF_ALL		: In   std_logic;
	     RAM_ADR_IS_AT_END_OFF_TEMPEXP	: In   std_logic;
	     RAM_ADR_IS_AT_END_OFF_MODUL	: In   std_logic;
	     RAM_ADR_IS_AT_END_OFF_PUBLICKEY	: In   std_logic;
	     RAM_ADR_IS_AT_END_OFF_PRIVATKEY	: In   std_logic;
	     RAM_ADR_IS_AT_END_OFF_ZERTPUB	: In   std_logic;
	     RAM_ADR_IS_AT_END_OFF_ZERTMODUL	: In   std_logic;
	     INVERT : out STD_LOGIC );

    end component;

    signal RAM_MODE				: STD_LOGIC_VECTOR(5 downto 0);
    signal RAM_ADR_I				: STD_LOGIC_VECTOR(7 downto 0);
    signal RAM_ADR_IS_AT_END_OFF_ALL		: STD_LOGIC;
    signal RAM_ADR_IS_AT_END_OFF_TEMPEXP	: STD_LOGIC;
    signal RAM_ADR_IS_AT_END_OFF_MODUL		: STD_LOGIC;
    signal RAM_ADR_IS_AT_END_OFF_PUBLICKEY	: STD_LOGIC;
    signal RAM_ADR_IS_AT_END_OFF_PRIVATKEY	: STD_LOGIC;
    signal RAM_ADR_IS_AT_END_OFF_ZERTPUB	: STD_LOGIC;
    signal RAM_ADR_IS_AT_END_OFF_ZERTMODUL	: STD_LOGIC;

    signal INVERT : STD_LOGIC;
    
begin
    RAM_ADR <= RAM_ADR_I;

    I_RAM_COUNTER : RAM_COUNTER
      Port Map ( RAM_ADR => RAM_ADR_I,
		 CLK => CLK,
		 RESET => RESET,
		 RAM_MODE => RAM_MODE,
		 RAM_ADR_IS_AT_END_OFF_ALL => RAM_ADR_IS_AT_END_OFF_ALL,
		 RAM_ADR_IS_AT_END_OFF_TEMPEXP => RAM_ADR_IS_AT_END_OFF_TEMPEXP,
		 RAM_ADR_IS_AT_END_OFF_MODUL => RAM_ADR_IS_AT_END_OFF_MODUL,
		 RAM_ADR_IS_AT_END_OFF_PRIVATKEY => RAM_ADR_IS_AT_END_OFF_PRIVATKEY,
		 RAM_ADR_IS_AT_END_OFF_PUBLICKEY => RAM_ADR_IS_AT_END_OFF_PUBLICKEY,
		 RAM_ADR_IS_AT_END_OFF_ZERTMODUL => RAM_ADR_IS_AT_END_OFF_ZERTMODUL,
		 RAM_ADR_IS_AT_END_OFF_ZERTPUB => RAM_ADR_IS_AT_END_OFF_ZERTPUB,
		 INVERT => INVERT);

    I_FSM_CORE : FSM_CORE
      Port map ( CARDCHANGE  => CARDCHANGE,
		 CLK => CLK,
		 CTRL => CTRL,
		 CTRL_CHANGE => CTRL_CHANGE,
		 DATA_VALID => DATA_VALID,
		 DES_BUFFER_FREE => DES_BUFFER_FREE,
		 DES_DATA_READY => DES_DATA_READY,
		 DES_ERR => DES_ERR,
		 DES_PARITY => DES_PARITY,
		 DOUT_EMPTY => DOUT_EMPTY,
		 EQUAL => EQUAL,
		 RESET => RESET,
		 RSA_NEXTEXP => RSA_NEXTEXP,
		 RSA_READY => RSA_READY,
		 BUSY => BUSY,
		 DES_BUFFER_FREE_SET => DES_BUFFER_FREE_SET,
		 DES_DATA_IS_KEY => DES_DATA_IS_KEY,
		 DES_DATA_READY_SET => DES_DATA_READY_SET,
		 DES_IN_EN => DES_IN_EN,
		 DES_MODE => DES_MODE,
		 DEST_REG => DEST_REG,
		 ENABLE_TEST => ENABLE_TEST,
		 EQ_REG => EQ_REG,
		 INT => INT,
		 RAM_SEL => RAM_SEL,
		 RSA_GO => RSA_GO,
		 RSA_SEL => RSA_SEL,
		 RSA_VAL_ACC => RSA_VAL_ACC,
		 SOURCE_REG => SOURCE_REG,
		 STATE_EN => STATE_EN,
		 STATUS => STATUS,
		 RAM_MODE => RAM_MODE,
		 RAM_ADR_IS_AT_END_OFF_ALL => RAM_ADR_IS_AT_END_OFF_ALL,
		 RAM_ADR_IS_AT_END_OFF_TEMPEXP => RAM_ADR_IS_AT_END_OFF_TEMPEXP,
		 RAM_ADR_IS_AT_END_OFF_MODUL => RAM_ADR_IS_AT_END_OFF_MODUL,
		 RAM_ADR_IS_AT_END_OFF_PRIVATKEY => RAM_ADR_IS_AT_END_OFF_PRIVATKEY,
		 RAM_ADR_IS_AT_END_OFF_PUBLICKEY => RAM_ADR_IS_AT_END_OFF_PUBLICKEY,
		 RAM_ADR_IS_AT_END_OFF_ZERTMODUL => RAM_ADR_IS_AT_END_OFF_ZERTMODUL,
		 RAM_ADR_IS_AT_END_OFF_ZERTPUB => RAM_ADR_IS_AT_END_OFF_ZERTPUB,
		 INVERT => INVERT );

end BEHAVIORAL;

