
----------------------------------------------------------------------------
--  This file is a part of the LEON VHDL model
--  Copyright (C) 1999  European Space Agency (ESA)
--
--  This library is free software; you can redistribute it and/or
--  modify it under the terms of the GNU Lesser General Public
--  License as published by the Free Software Foundation; either
--  version 2 of the License, or (at your option) any later version.
--
--  See the file COPYING.LGPL for the full details of the license.


-----------------------------------------------------------------------------
-- Entity: 	rstgen
-- File:	rstgen.vhd
-- Author:	Jiri Gaisler - ESA/ESTEC
-- Description:	Internal reset is generated by this unit.

------------------------------------------------------------------------------
-- Version control:
-- 11-10-1998:	First implemetation
-- 26-09-1999:	Release 1.0
-- 08-12-1999:	Asynchronous clear of reset registers
------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use work.config.all;
use work.iface.all;

entity rstgen is
port (
    resetn : in  std_logic;
    pcirst : in  std_logic;
    clk    : in  clk_type;
    rst    : out rst_type
);
end;

architecture rtl of rstgen is
signal rstr, rstrin : std_logic_vector(3 downto 0);
signal rstall : std_logic;

begin

-- reset generation

  rstall <= resetn and pcirst when PCIEN else resetn;


  reg1 : process (clk,rstall) begin
    if rstall = '0' then rstr <= "0000";
    elsif rising_edge(clk) then rstr <= rstr(2 downto 0) & '1'; end if;
  end process;

  rst.syncrst <= rstr(3);
  rst.rawrst  <= rstall;

end;

