-------------------------------------------------------------------------------
-- Crypto Chip
-- Copyright (C) 1999, Projektgruppe WS98/99
-- University of Stuttgart / Department of Computer Science / IFI-RA
-------------------------------------------------------------------------------
-- Designers:        Joerg Holzhauer
-- Group    :        DES
-------------------------------------------------------------------------------
-- Design Unit Name: DES_S7_Box
-- Purpose:          Gate for the DES-module-core for the cryptochip "pg99"
--
-- File Name:        s7.vhd
-------------------------------------------------------------------------------
-- Simulator :       SYNOPSIS VHDL System Simulator (VSS) Version 3.2.a
-------------------------------------------------------------------------------
-- Date    09.11.98 |  Changes
--                  |
--                  |
-------------------------------------------------------------------------------

-------------------------------------------------------------------------------
-- contents :        port- and behaviour-description of
--                   one Gate of the DES-Module
--
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;
entity DES_S7_Box is
  port (i :in STD_LOGIC_VECTOR(0 to 5);
        o :out STD_LOGIC_VECTOR(0 to 3));
end DES_S7_Box;

architecture behavorial of DES_S7_Box is
begin
with i select
o(0) <= '1' when "000010"|
"000110"|
"001000"|
"001100"|
"001110"|
"010010"|
"010100"|
"011010"|
"000001"|
"000101"|
"001011"|
"001111"|
"010001"|
"010111"|
"011011"|
"011101"|
"100100"|
"100110"|
"101000"|
"101110"|
"110000"|
"110010"|
"110110"|
"111100"|
"100011"|
"100101"|
"100111"|
"101101"|
"110001"|
"110111"|
"111001"|
"111111",
'0' when others;
with i select
o(1) <= '1' when "000000"|
"000110"|
"001000"|
"001110"|
"010010"|
"010110"|
"011000"|
"011100"|
"000001"|
"000111"|
"001001"|
"010001"|
"010101"|
"010111"|
"011011"|
"011111"|
"100010"|
"100110"|
"101000"|
"101100"|
"101110"|
"110010"|
"110100"|
"111010"|
"100001"|
"100101"|
"101011"|
"101111"|
"110011"|
"110111"|
"111001"|
"111111",
'0' when others;
with i select
o(2) <= '1' when "000010"|
"000100"|
"000110"|
"001000"|
"010000"|
"010110"|
"011010"|
"011100"|
"000101"|
"000111"|
"001111"|
"010001"|
"010011"|
"011001"|
"011011"|
"011111"|
"100100"|
"101010"|
"101100"|
"101110"|
"110000"|
"110010"|
"110100"|
"111110"|
"100001"|
"100011"|
"101101"|
"101111"|
"110111"|
"111001"|
"111011"|
"111101",
'0' when others;
with i select
o(3) <= '1' when "000010"|
"001000"|
"001110"|
"010000"|
"010100"|
"010110"|
"011000"|
"011110"|
"000001"|
"000101"|
"000111"|
"001011"|
"001101"|
"010011"|
"010101"|
"011011"|
"100000"|
"100100"|
"100110"|
"101010"|
"101100"|
"110010"|
"111010"|
"111100"|
"100011"|
"100101"|
"101001"|
"101111"|
"110001"|
"110011"|
"110111"|
"111101",
'0' when others;
end behavorial;
